module decoder_90836_06260 (
	debug_req_i,
	pc_i,
	is_compressed_i,
	compressed_instr_i,
	is_illegal_i,
	instruction_i,
	is_macro_instr_i,
	is_last_macro_instr_i,
	is_double_rd_macro_instr_i,
	branch_predict_i,
	ex_i,
	irq_i,
	irq_ctrl_i,
	priv_lvl_i,
	v_i,
	debug_mode_i,
	fs_i,
	vfs_i,
	frm_i,
	vs_i,
	tvm_i,
	tw_i,
	vtw_i,
	tsr_i,
	hu_i,
	instruction_o,
	orig_instr_o,
	is_control_flow_instr_o
);
	// removed localparam type branchpredict_sbe_t_branchpredict_sbe_t_CVA6Cfg_type
	parameter [17102:0] branchpredict_sbe_t_branchpredict_sbe_t_CVA6Cfg = 0;
	// removed localparam type exception_t_exception_t_CVA6Cfg_type
	parameter [17102:0] exception_t_exception_t_CVA6Cfg = 0;
	// removed localparam type interrupts_t_interrupts_t_CVA6Cfg_type
	parameter [17102:0] interrupts_t_interrupts_t_CVA6Cfg = 0;
	// removed localparam type irq_ctrl_t_irq_ctrl_t_CVA6Cfg_type
	parameter [17102:0] irq_ctrl_t_irq_ctrl_t_CVA6Cfg = 0;
	// removed localparam type scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg_type
	parameter [17102:0] scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg = 0;
	reg _sv2v_0;
	// removed import ariane_pkg::*;
	// Trace: core/decoder.sv:25:15
	localparam config_pkg_NrMaxRules = 16;
	// removed localparam type config_pkg_cache_type_t
	// removed localparam type config_pkg_noc_type_e
	// removed localparam type config_pkg_vm_mode_t
	// removed localparam type config_pkg_cva6_cfg_t
	localparam [17102:0] config_pkg_cva6_cfg_empty = 17103'd0;
	parameter [17102:0] CVA6Cfg = config_pkg_cva6_cfg_empty;
	// Trace: core/decoder.sv:26:20
	// removed localparam type branchpredict_sbe_t
	// Trace: core/decoder.sv:27:20
	// removed localparam type exception_t
	// Trace: core/decoder.sv:28:20
	// removed localparam type irq_ctrl_t
	// Trace: core/decoder.sv:29:20
	// removed localparam type scoreboard_entry_t
	// Trace: core/decoder.sv:30:20
	// removed localparam type interrupts_t
	// Trace: core/decoder.sv:31:15
	parameter [(((((((((interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + interrupts_t_interrupts_t_CVA6Cfg[17102-:32]) + interrupts_t_interrupts_t_CVA6Cfg[17102-:32]) + interrupts_t_interrupts_t_CVA6Cfg[17102-:32]) + interrupts_t_interrupts_t_CVA6Cfg[17102-:32]) + interrupts_t_interrupts_t_CVA6Cfg[17102-:32]) + interrupts_t_interrupts_t_CVA6Cfg[17102-:32]) + interrupts_t_interrupts_t_CVA6Cfg[17102-:32]) + interrupts_t_interrupts_t_CVA6Cfg[17102-:32]) + interrupts_t_interrupts_t_CVA6Cfg[17102-:32]) - 1:0] INTERRUPTS = 1'sb0;
	// Trace: core/decoder.sv:34:5
	input wire debug_req_i;
	// Trace: core/decoder.sv:36:5
	input wire [CVA6Cfg[17070-:32] - 1:0] pc_i;
	// Trace: core/decoder.sv:38:5
	input wire is_compressed_i;
	// Trace: core/decoder.sv:40:5
	input wire [15:0] compressed_instr_i;
	// Trace: core/decoder.sv:42:5
	input wire is_illegal_i;
	// Trace: core/decoder.sv:44:5
	input wire [31:0] instruction_i;
	// Trace: core/decoder.sv:46:5
	input wire is_macro_instr_i;
	// Trace: core/decoder.sv:48:5
	input wire is_last_macro_instr_i;
	// Trace: core/decoder.sv:50:5
	input wire is_double_rd_macro_instr_i;
	// Trace: core/decoder.sv:52:5
	input wire [(3 + branchpredict_sbe_t_branchpredict_sbe_t_CVA6Cfg[17070-:32]) - 1:0] branch_predict_i;
	// Trace: core/decoder.sv:54:5
	input wire [((exception_t_exception_t_CVA6Cfg[17102-:32] + exception_t_exception_t_CVA6Cfg[17102-:32]) + exception_t_exception_t_CVA6Cfg[17006-:32]) + 33:0] ex_i;
	// Trace: core/decoder.sv:56:5
	input wire [1:0] irq_i;
	// Trace: core/decoder.sv:58:5
	input wire [(((irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32]) + irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32]) + irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32]) + 1:0] irq_ctrl_i;
	// Trace: core/decoder.sv:60:5
	// removed localparam type riscv_priv_lvl_t
	input wire [1:0] priv_lvl_i;
	// Trace: core/decoder.sv:62:5
	input wire v_i;
	// Trace: core/decoder.sv:64:5
	input wire debug_mode_i;
	// Trace: core/decoder.sv:66:5
	// removed localparam type riscv_xs_t
	input wire [1:0] fs_i;
	// Trace: core/decoder.sv:68:5
	input wire [1:0] vfs_i;
	// Trace: core/decoder.sv:70:5
	input wire [2:0] frm_i;
	// Trace: core/decoder.sv:72:5
	input wire [1:0] vs_i;
	// Trace: core/decoder.sv:74:5
	input wire tvm_i;
	// Trace: core/decoder.sv:76:5
	input wire tw_i;
	// Trace: core/decoder.sv:78:5
	input wire vtw_i;
	// Trace: core/decoder.sv:80:5
	input wire tsr_i;
	// Trace: core/decoder.sv:82:5
	input wire hu_i;
	// Trace: core/decoder.sv:84:5
	output reg [((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4:0] instruction_o;
	// Trace: core/decoder.sv:86:5
	output reg [31:0] orig_instr_o;
	// Trace: core/decoder.sv:88:5
	output reg is_control_flow_instr_o;
	// Trace: core/decoder.sv:90:3
	reg illegal_instr;
	// Trace: core/decoder.sv:91:3
	reg illegal_instr_bm;
	// Trace: core/decoder.sv:92:3
	reg illegal_instr_zic;
	// Trace: core/decoder.sv:93:3
	reg illegal_instr_non_bm;
	// Trace: core/decoder.sv:94:3
	reg virtual_illegal_instr;
	// Trace: core/decoder.sv:96:3
	reg ecall;
	// Trace: core/decoder.sv:98:3
	reg ebreak;
	// Trace: core/decoder.sv:100:3
	reg check_fprm;
	// Trace: core/decoder.sv:101:3
	// removed localparam type riscv_atype_t
	// removed localparam type riscv_itype_t
	// removed localparam type riscv_r4type_t
	// removed localparam type riscv_rftype_t
	// removed localparam type riscv_rtype_t
	// removed localparam type riscv_rvftype_t
	// removed localparam type riscv_stype_t
	// removed localparam type riscv_utype_t
	// removed localparam type riscv_instruction_t
	wire [31:0] instr;
	// Trace: core/decoder.sv:102:3
	assign instr = instruction_i;
	// Trace: core/decoder.sv:104:3
	reg [31:0] tinst;
	// Trace: core/decoder.sv:108:3
	reg [3:0] imm_select;
	// Trace: core/decoder.sv:119:3
	reg [CVA6Cfg[17102-:32] - 1:0] imm_i_type;
	// Trace: core/decoder.sv:120:3
	reg [CVA6Cfg[17102-:32] - 1:0] imm_s_type;
	// Trace: core/decoder.sv:121:3
	reg [CVA6Cfg[17102-:32] - 1:0] imm_sb_type;
	// Trace: core/decoder.sv:122:3
	reg [CVA6Cfg[17102-:32] - 1:0] imm_u_type;
	// Trace: core/decoder.sv:123:3
	reg [CVA6Cfg[17102-:32] - 1:0] imm_uj_type;
	// Trace: core/decoder.sv:124:3
	reg [CVA6Cfg[17102-:32] - 1:0] imm_bi_type;
	// Trace: core/decoder.sv:129:3
	wire is_accel;
	// Trace: core/decoder.sv:130:3
	wire [((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4:0] acc_instruction;
	// Trace: core/decoder.sv:131:3
	wire acc_illegal_instr;
	// Trace: core/decoder.sv:132:3
	wire acc_is_control_flow_instr;
	// Trace: core/decoder.sv:134:3
	generate
		if (CVA6Cfg[16369]) begin : gen_accel_decoder
			// Trace: core/decoder.sv:138:5
			cva6_accel_first_pass_decoder_AA251_75519 #(
				.scoreboard_entry_t_scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg(scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg),
				.CVA6Cfg(CVA6Cfg)
			) i_accel_decoder(
				.instruction_i(instruction_i),
				.fs_i(fs_i),
				.vs_i(vs_i),
				.is_accel_o(is_accel),
				.instruction_o(acc_instruction),
				.illegal_instr_o(acc_illegal_instr),
				.is_control_flow_instr_o(acc_is_control_flow_instr)
			);
		end
		else begin : genblk1
			// Trace: core/decoder.sv:152:5
			assign is_accel = 1'b0;
			// Trace: core/decoder.sv:153:5
			assign acc_instruction = 1'sb0;
			// Trace: core/decoder.sv:154:5
			assign acc_illegal_instr = 1'b1;
			// Trace: core/decoder.sv:155:5
			assign acc_is_control_flow_instr = 1'b0;
		end
	endgenerate
	// Trace: core/decoder.sv:158:3
	// removed localparam type ariane_pkg_fu_op
	// removed localparam type ariane_pkg_fu_t
	localparam riscv_OpcodeAmo = 7'b0101111;
	localparam riscv_OpcodeAuipc = 7'b0010111;
	localparam riscv_OpcodeBranch = 7'b1100011;
	localparam riscv_OpcodeJal = 7'b1101111;
	localparam riscv_OpcodeJalr = 7'b1100111;
	localparam riscv_OpcodeLoad = 7'b0000011;
	localparam riscv_OpcodeLoadFp = 7'b0000111;
	localparam riscv_OpcodeLui = 7'b0110111;
	localparam riscv_OpcodeMadd = 7'b1000011;
	localparam riscv_OpcodeMiscMem = 7'b0001111;
	localparam riscv_OpcodeMsub = 7'b1000111;
	localparam riscv_OpcodeNmadd = 7'b1001111;
	localparam riscv_OpcodeNmsub = 7'b1001011;
	localparam riscv_OpcodeOp = 7'b0110011;
	localparam riscv_OpcodeOp32 = 7'b0111011;
	localparam riscv_OpcodeOpFp = 7'b1010011;
	localparam riscv_OpcodeOpImm = 7'b0010011;
	localparam riscv_OpcodeOpImm32 = 7'b0011011;
	localparam riscv_OpcodeStore = 7'b0100011;
	localparam riscv_OpcodeStoreFp = 7'b0100111;
	localparam riscv_OpcodeSystem = 7'b1110011;
	always @(*) begin : decoder
		if (_sv2v_0)
			;
		// Trace: core/decoder.sv:160:5
		imm_select = 4'd0;
		// Trace: core/decoder.sv:161:5
		is_control_flow_instr_o = 1'b0;
		// Trace: core/decoder.sv:162:5
		illegal_instr = 1'b0;
		// Trace: core/decoder.sv:163:5
		illegal_instr_non_bm = 1'b0;
		// Trace: core/decoder.sv:164:5
		illegal_instr_bm = 1'b0;
		// Trace: core/decoder.sv:165:5
		illegal_instr_zic = 1'b0;
		// Trace: core/decoder.sv:166:5
		virtual_illegal_instr = 1'b0;
		// Trace: core/decoder.sv:167:5
		instruction_o[scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))-:((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))))) + 1)] = pc_i;
		// Trace: core/decoder.sv:168:5
		instruction_o[scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))-:((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) >= (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + 1)] = 1'sb0;
		// Trace: core/decoder.sv:169:5
		instruction_o[27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 4'd0;
		// Trace: core/decoder.sv:170:5
		instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd0;
		// Trace: core/decoder.sv:171:5
		instruction_o[15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 1'sb0;
		// Trace: core/decoder.sv:172:5
		instruction_o[10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 1'sb0;
		// Trace: core/decoder.sv:173:5
		instruction_o[5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 1'sb0;
		// Trace: core/decoder.sv:174:5
		instruction_o[1 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))] = 1'b0;
		// Trace: core/decoder.sv:175:5
		instruction_o[4] = is_compressed_i;
		// Trace: core/decoder.sv:176:5
		instruction_o[3] = is_macro_instr_i;
		// Trace: core/decoder.sv:177:5
		instruction_o[2] = is_last_macro_instr_i;
		// Trace: core/decoder.sv:178:5
		instruction_o[1] = is_double_rd_macro_instr_i;
		// Trace: core/decoder.sv:179:5
		instruction_o[2 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))] = 1'b0;
		// Trace: core/decoder.sv:180:5
		instruction_o[(3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4-:(((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4) >= 5 ? (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 0 : 6 - ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))] = branch_predict_i;
		// Trace: core/decoder.sv:181:5
		instruction_o[0] = 1'b0;
		// Trace: core/decoder.sv:182:5
		tinst = 1'sb0;
		// Trace: core/decoder.sv:183:5
		ecall = 1'b0;
		// Trace: core/decoder.sv:184:5
		ebreak = 1'b0;
		// Trace: core/decoder.sv:185:5
		check_fprm = 1'b0;
		// Trace: core/decoder.sv:187:5
		if (~ex_i[0])
			// Trace: core/decoder.sv:188:7
			case (instr[6-:7])
				riscv_OpcodeSystem: begin
					// Trace: core/decoder.sv:190:11
					instruction_o[27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 4'd6;
					// Trace: core/decoder.sv:191:11
					instruction_o[15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[19-:5];
					// Trace: core/decoder.sv:192:11
					instruction_o[10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[24-:5];
					// Trace: core/decoder.sv:193:11
					instruction_o[5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[11-:5];
					// Trace: core/decoder.sv:195:11
					(* full_case, parallel_case *)
					case (instr[14-:3])
						3'b000: begin
							// Trace: core/decoder.sv:198:15
							if ((instr[19-:5] != {5 {1'sb0}}) || (instr[11-:5] != {5 {1'sb0}})) begin
								begin
									// Trace: core/decoder.sv:199:17
									if (CVA6Cfg[16543] && v_i)
										// Trace: core/decoder.sv:200:19
										virtual_illegal_instr = 1'b1;
									else
										// Trace: core/decoder.sv:202:19
										illegal_instr = 1'b1;
								end
							end
							case (instr[31-:12])
								12'b000000000000:
									// Trace: core/decoder.sv:208:24
									ecall = 1'b1;
								12'b000000000001:
									// Trace: core/decoder.sv:210:24
									ebreak = 1'b1;
								12'b000100000010:
									// Trace: core/decoder.sv:213:19
									if (CVA6Cfg[16366]) begin
										// Trace: core/decoder.sv:214:21
										instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd24;
										// Trace: core/decoder.sv:217:21
										if (CVA6Cfg[16365] && (priv_lvl_i == 2'b00)) begin
											// Trace: core/decoder.sv:218:23
											if (CVA6Cfg[16543] && v_i)
												// Trace: core/decoder.sv:219:25
												virtual_illegal_instr = 1'b1;
											else
												// Trace: core/decoder.sv:221:25
												illegal_instr = 1'b1;
											// Trace: core/decoder.sv:224:23
											instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd0;
										end
										if ((priv_lvl_i == 2'b01) && tsr_i) begin
											// Trace: core/decoder.sv:228:23
											if (CVA6Cfg[16543] && v_i)
												// Trace: core/decoder.sv:229:25
												virtual_illegal_instr = 1'b1;
											else
												// Trace: core/decoder.sv:231:25
												illegal_instr = 1'b1;
											// Trace: core/decoder.sv:234:23
											instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd0;
										end
									end
									else begin
										// Trace: core/decoder.sv:237:21
										illegal_instr = 1'b1;
										// Trace: core/decoder.sv:238:21
										instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd0;
									end
								12'b001100000010: begin
									// Trace: core/decoder.sv:243:19
									instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd23;
									// Trace: core/decoder.sv:246:19
									if ((CVA6Cfg[16366] && (priv_lvl_i == 2'b01)) || (CVA6Cfg[16365] && (priv_lvl_i == 2'b00)))
										// Trace: core/decoder.sv:247:21
										illegal_instr = 1'b1;
								end
								12'b011110110010: begin
									// Trace: core/decoder.sv:251:19
									instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd25;
									// Trace: core/decoder.sv:252:19
									if (CVA6Cfg[1321])
										// Trace: core/decoder.sv:254:21
										illegal_instr = (!debug_mode_i ? 1'b1 : illegal_instr);
									else
										// Trace: core/decoder.sv:256:21
										illegal_instr = 1'b1;
								end
								12'b000100000101: begin
									// Trace: core/decoder.sv:261:19
									instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd27;
									// Trace: core/decoder.sv:264:19
									if ((CVA6Cfg[16366] && (priv_lvl_i == 2'b01)) && tw_i) begin
										// Trace: core/decoder.sv:265:21
										illegal_instr = 1'b1;
										// Trace: core/decoder.sv:266:21
										instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd0;
									end
									if ((((CVA6Cfg[16543] && (priv_lvl_i == 2'b01)) && v_i) && vtw_i) && !tw_i) begin
										// Trace: core/decoder.sv:269:21
										virtual_illegal_instr = 1'b1;
										// Trace: core/decoder.sv:270:21
										instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd0;
									end
									if (CVA6Cfg[16365] && (priv_lvl_i == 2'b00)) begin
										// Trace: core/decoder.sv:274:21
										if (CVA6Cfg[16543] && v_i)
											// Trace: core/decoder.sv:274:45
											virtual_illegal_instr = 1'b1;
										else
											// Trace: core/decoder.sv:275:26
											illegal_instr = 1'b1;
										// Trace: core/decoder.sv:276:21
										instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd0;
									end
								end
								default:
									// Trace: core/decoder.sv:281:19
									if (instr[31:25] == 7'b0001001) begin
										// Trace: core/decoder.sv:285:21
										if (CVA6Cfg[16543] && v_i)
											// Trace: core/decoder.sv:286:23
											virtual_illegal_instr = (priv_lvl_i == 2'b01 ? 1'b0 : 1'b1);
										else
											// Trace: core/decoder.sv:288:23
											illegal_instr = ((CVA6Cfg[16366] && |{priv_lvl_i == 2'b11, priv_lvl_i == 2'b01}) && (instr[11-:5] == {5 {1'sb0}}) ? 1'b0 : 1'b1);
										// Trace: core/decoder.sv:290:21
										instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd30;
										if ((CVA6Cfg[16366] && (priv_lvl_i == 2'b01)) && tvm_i) begin
											begin
												// Trace: core/decoder.sv:293:23
												if (CVA6Cfg[16543] && v_i)
													// Trace: core/decoder.sv:293:47
													virtual_illegal_instr = 1'b1;
												else
													// Trace: core/decoder.sv:294:28
													illegal_instr = 1'b1;
											end
										end
									end
									else if (CVA6Cfg[16543]) begin
										begin
											// Trace: core/decoder.sv:297:21
											if (instr[31:25] == 7'b0010001) begin
												// Trace: core/decoder.sv:300:23
												if (v_i)
													// Trace: core/decoder.sv:301:25
													virtual_illegal_instr = 1'b1;
												else
													// Trace: core/decoder.sv:303:25
													illegal_instr = (|{priv_lvl_i == 2'b11, priv_lvl_i == 2'b01} ? 1'b0 : 1'b1);
												// Trace: core/decoder.sv:305:23
												instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd31;
											end
											else if (instr[31:25] == 7'b0110001) begin
												// Trace: core/decoder.sv:309:23
												if (v_i)
													// Trace: core/decoder.sv:310:25
													virtual_illegal_instr = 1'b1;
												else
													// Trace: core/decoder.sv:312:25
													illegal_instr = (|{priv_lvl_i == 2'b11, priv_lvl_i == 2'b01} ? 1'b0 : 1'b1);
												// Trace: core/decoder.sv:314:23
												instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd32;
												if (((priv_lvl_i == 2'b01) && !v_i) && tvm_i)
													// Trace: core/decoder.sv:316:77
													illegal_instr = 1'b1;
											end
											else
												// Trace: core/decoder.sv:318:23
												illegal_instr = 1'b1;
										end
									end
									else
										// Trace: core/decoder.sv:321:21
										illegal_instr = 1'b1;
							endcase
						end
						3'b100:
							// Trace: core/decoder.sv:328:15
							if (CVA6Cfg[16543]) begin
								// Trace: core/decoder.sv:329:17
								if (instr[25] != 1'b0) begin
									// Trace: core/decoder.sv:330:19
									instruction_o[27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 4'd2;
									// Trace: core/decoder.sv:331:19
									imm_select = 4'd0;
									// Trace: core/decoder.sv:332:19
									instruction_o[15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[19-:5];
									// Trace: core/decoder.sv:333:19
									instruction_o[10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[24-:5];
								end
								else begin
									// Trace: core/decoder.sv:335:19
									instruction_o[27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 4'd1;
									// Trace: core/decoder.sv:336:19
									imm_select = 4'd0;
									// Trace: core/decoder.sv:337:19
									instruction_o[15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[19-:5];
									// Trace: core/decoder.sv:338:19
									instruction_o[5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[11-:5];
								end
								if (v_i)
									// Trace: core/decoder.sv:342:26
									virtual_illegal_instr = 1'b1;
								else if (!hu_i && (priv_lvl_i == 2'b00))
									// Trace: core/decoder.sv:344:68
									illegal_instr = 1'b1;
								(* full_case, parallel_case *)
								case (instr[31-:7])
									7'b0110000: begin
										// Trace: core/decoder.sv:347:21
										if (instr[24-:5] == 5'b00000)
											// Trace: core/decoder.sv:348:23
											instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd48;
										if (instr[24-:5] == 5'b00001)
											// Trace: core/decoder.sv:351:23
											instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd49;
									end
									7'b0110010: begin
										// Trace: core/decoder.sv:355:21
										if (instr[24-:5] == 5'b00000)
											// Trace: core/decoder.sv:356:23
											instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd50;
										if (instr[24-:5] == 5'b00001)
											// Trace: core/decoder.sv:359:23
											instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd51;
										if (instr[24-:5] == 5'b00011)
											// Trace: core/decoder.sv:362:23
											instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd52;
									end
									7'b0110100: begin
										// Trace: core/decoder.sv:366:21
										if (instr[24-:5] == 5'b00000)
											// Trace: core/decoder.sv:367:23
											instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd53;
										if (instr[24-:5] == 5'b00001)
											// Trace: core/decoder.sv:370:23
											instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd58;
										if (instr[24-:5] == 5'b00011)
											// Trace: core/decoder.sv:373:23
											instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd54;
									end
									7'b0110001:
										// Trace: core/decoder.sv:376:32
										instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd55;
									7'b0110011:
										// Trace: core/decoder.sv:377:32
										instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd56;
									7'b0110101:
										// Trace: core/decoder.sv:378:32
										instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd57;
									7'b0110110:
										// Trace: core/decoder.sv:379:32
										instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd59;
									7'b0110111:
										// Trace: core/decoder.sv:380:32
										instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd60;
									default:
										// Trace: core/decoder.sv:381:28
										illegal_instr = 1'b1;
								endcase
								// Trace: core/decoder.sv:384:17
								tinst = {instr[31-:7], instr[24-:5], 5'b00000, instr[14-:3], instr[11-:5], instr[6-:7]};
							end
							else
								// Trace: core/decoder.sv:393:17
								illegal_instr = 1'b1;
						3'b001: begin
							// Trace: core/decoder.sv:398:15
							imm_select = 4'd1;
							// Trace: core/decoder.sv:399:15
							instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd33;
						end
						3'b010: begin
							// Trace: core/decoder.sv:403:15
							imm_select = 4'd1;
							// Trace: core/decoder.sv:405:15
							if (instr[19-:5] == 5'b00000)
								// Trace: core/decoder.sv:405:44
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd34;
							else
								// Trace: core/decoder.sv:406:20
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd35;
						end
						3'b011: begin
							// Trace: core/decoder.sv:410:15
							imm_select = 4'd1;
							// Trace: core/decoder.sv:412:15
							if (instr[19-:5] == 5'b00000)
								// Trace: core/decoder.sv:412:44
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd34;
							else
								// Trace: core/decoder.sv:413:20
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd36;
						end
						3'b101: begin
							// Trace: core/decoder.sv:417:15
							instruction_o[15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[19-:5];
							// Trace: core/decoder.sv:418:15
							imm_select = 4'd1;
							// Trace: core/decoder.sv:419:15
							instruction_o[2 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))] = 1'b1;
							// Trace: core/decoder.sv:420:15
							instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd33;
						end
						3'b110: begin
							// Trace: core/decoder.sv:423:15
							instruction_o[15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[19-:5];
							// Trace: core/decoder.sv:424:15
							imm_select = 4'd1;
							// Trace: core/decoder.sv:425:15
							instruction_o[2 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))] = 1'b1;
							// Trace: core/decoder.sv:427:15
							if (instr[19-:5] == 5'b00000)
								// Trace: core/decoder.sv:427:44
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd34;
							else
								// Trace: core/decoder.sv:428:20
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd35;
						end
						3'b111: begin
							// Trace: core/decoder.sv:431:15
							instruction_o[15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[19-:5];
							// Trace: core/decoder.sv:432:15
							imm_select = 4'd1;
							// Trace: core/decoder.sv:433:15
							instruction_o[2 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))] = 1'b1;
							// Trace: core/decoder.sv:435:15
							if (instr[19-:5] == 5'b00000)
								// Trace: core/decoder.sv:435:44
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd34;
							else
								// Trace: core/decoder.sv:436:20
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd36;
						end
						default:
							// Trace: core/decoder.sv:438:22
							illegal_instr = 1'b1;
					endcase
				end
				riscv_OpcodeMiscMem: begin
					// Trace: core/decoder.sv:443:11
					instruction_o[27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 4'd6;
					// Trace: core/decoder.sv:444:11
					instruction_o[15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 1'sb0;
					// Trace: core/decoder.sv:445:11
					instruction_o[10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 1'sb0;
					// Trace: core/decoder.sv:446:11
					instruction_o[5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 1'sb0;
					// Trace: core/decoder.sv:448:11
					case (instr[14-:3])
						3'b000:
							// Trace: core/decoder.sv:451:21
							instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd28;
						3'b001:
							// Trace: core/decoder.sv:453:21
							instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd29;
						default:
							// Trace: core/decoder.sv:455:22
							illegal_instr = 1'b1;
					endcase
				end
				riscv_OpcodeOp:
					// Trace: core/decoder.sv:466:11
					if (instr[31-:2] == 2'b10) begin
						begin
							// Trace: core/decoder.sv:468:13
							if (((CVA6Cfg[16471] && CVA6Cfg[16540]) && (fs_i != 2'b00)) && ((CVA6Cfg[16543] && (!v_i || (vfs_i != 2'b00))) || !CVA6Cfg[16543])) begin : sv2v_autoblock_1
								// Trace: core/decoder.sv:469:15
								reg allow_replication;
								// Trace: core/decoder.sv:471:15
								instruction_o[27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 4'd8;
								// Trace: core/decoder.sv:472:15
								instruction_o[15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[19-:5];
								// Trace: core/decoder.sv:473:15
								instruction_o[10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[24-:5];
								// Trace: core/decoder.sv:474:15
								instruction_o[5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[11-:5];
								// Trace: core/decoder.sv:475:15
								check_fprm = 1'b1;
								// Trace: core/decoder.sv:476:15
								allow_replication = 1'b1;
								// Trace: core/decoder.sv:478:15
								(* full_case, parallel_case *)
								case (instr[29-:5])
									5'b00001: begin
										// Trace: core/decoder.sv:480:19
										instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd104;
										// Trace: core/decoder.sv:481:19
										instruction_o[15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 1'sb0;
										// Trace: core/decoder.sv:482:19
										instruction_o[10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[19-:5];
										// Trace: core/decoder.sv:483:19
										imm_select = 4'd1;
									end
									5'b00010: begin
										// Trace: core/decoder.sv:486:19
										instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd105;
										// Trace: core/decoder.sv:487:19
										instruction_o[15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 1'sb0;
										// Trace: core/decoder.sv:488:19
										instruction_o[10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[19-:5];
										// Trace: core/decoder.sv:489:19
										imm_select = 4'd1;
									end
									5'b00011:
										// Trace: core/decoder.sv:492:17
										instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd106;
									5'b00100:
										// Trace: core/decoder.sv:494:17
										instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd107;
									5'b00101: begin
										// Trace: core/decoder.sv:496:19
										instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd122;
										// Trace: core/decoder.sv:497:19
										check_fprm = 1'b0;
									end
									5'b00110: begin
										// Trace: core/decoder.sv:500:19
										instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd123;
										// Trace: core/decoder.sv:501:19
										check_fprm = 1'b0;
									end
									5'b00111: begin
										// Trace: core/decoder.sv:504:19
										instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd109;
										// Trace: core/decoder.sv:505:19
										allow_replication = 1'b0;
										// Trace: core/decoder.sv:506:19
										if (instr[24-:5] != 5'b00000)
											// Trace: core/decoder.sv:506:54
											illegal_instr = 1'b1;
									end
									5'b01000: begin
										// Trace: core/decoder.sv:509:19
										instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd110;
										// Trace: core/decoder.sv:510:19
										imm_select = 4'd2;
									end
									5'b01001: begin
										// Trace: core/decoder.sv:513:19
										instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd111;
										// Trace: core/decoder.sv:514:19
										imm_select = 4'd2;
									end
									5'b01100:
										// Trace: core/decoder.sv:517:19
										(* full_case, parallel_case *)
										if (instr[24-:5] == 5'b00000) begin
											// Trace: core/decoder.sv:519:23
											instruction_o[10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[19-:5];
											// Trace: core/decoder.sv:520:23
											if (instr[14])
												// Trace: core/decoder.sv:521:25
												instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd119;
											else
												// Trace: core/decoder.sv:522:28
												instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd118;
											// Trace: core/decoder.sv:523:23
											check_fprm = 1'b0;
										end
										else if (instr[24-:5] == 5'b00001) begin
											// Trace: core/decoder.sv:526:23
											instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd121;
											// Trace: core/decoder.sv:527:23
											check_fprm = 1'b0;
											// Trace: core/decoder.sv:528:23
											allow_replication = 1'b0;
										end
										else if (instr[24-:5] == 5'b00010)
											// Trace: core/decoder.sv:531:21
											instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd114;
										else if (instr[24-:5] == 5'b00011)
											// Trace: core/decoder.sv:533:21
											instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd115;
										else if ((instr[24-:5] | 5'b00011) == 5'b00111) begin
											// Trace: core/decoder.sv:535:23
											instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd116;
											// Trace: core/decoder.sv:536:23
											instruction_o[10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[11-:5];
											// Trace: core/decoder.sv:537:23
											imm_select = 4'd1;
											// Trace: core/decoder.sv:540:23
											(* full_case, parallel_case *)
											case (instr[21:20])
												2'b00:
													if (~CVA6Cfg[16437])
														// Trace: core/decoder.sv:542:55
														illegal_instr = 1'b1;
												2'b01:
													if (~CVA6Cfg[16435])
														// Trace: core/decoder.sv:543:59
														illegal_instr = 1'b1;
												2'b10:
													if (~CVA6Cfg[16436])
														// Trace: core/decoder.sv:544:56
														illegal_instr = 1'b1;
												2'b11:
													if (~CVA6Cfg[16434])
														// Trace: core/decoder.sv:545:55
														illegal_instr = 1'b1;
												default:
													// Trace: core/decoder.sv:546:34
													illegal_instr = 1'b1;
											endcase
										end
										else
											// Trace: core/decoder.sv:549:30
											illegal_instr = 1'b1;
									5'b01101: begin
										// Trace: core/decoder.sv:553:19
										check_fprm = 1'b0;
										// Trace: core/decoder.sv:554:19
										instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd124;
									end
									5'b01110: begin
										// Trace: core/decoder.sv:557:19
										check_fprm = 1'b0;
										// Trace: core/decoder.sv:558:19
										instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd125;
									end
									5'b01111: begin
										// Trace: core/decoder.sv:561:19
										check_fprm = 1'b0;
										// Trace: core/decoder.sv:562:19
										instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd126;
									end
									5'b10000: begin
										// Trace: core/decoder.sv:565:19
										check_fprm = 1'b0;
										// Trace: core/decoder.sv:566:19
										instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd127;
									end
									5'b10001: begin
										// Trace: core/decoder.sv:569:19
										check_fprm = 1'b0;
										// Trace: core/decoder.sv:570:19
										instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd128;
									end
									5'b10010: begin
										// Trace: core/decoder.sv:573:19
										check_fprm = 1'b0;
										// Trace: core/decoder.sv:574:19
										instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd129;
									end
									5'b10011: begin
										// Trace: core/decoder.sv:577:19
										check_fprm = 1'b0;
										// Trace: core/decoder.sv:578:19
										instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd130;
									end
									5'b10100: begin
										// Trace: core/decoder.sv:581:19
										check_fprm = 1'b0;
										// Trace: core/decoder.sv:582:19
										instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd131;
									end
									5'b10101: begin
										// Trace: core/decoder.sv:585:19
										check_fprm = 1'b0;
										// Trace: core/decoder.sv:586:19
										instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd132;
									end
									5'b11000: begin
										// Trace: core/decoder.sv:589:19
										instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd133;
										// Trace: core/decoder.sv:590:19
										imm_select = 4'd2;
										// Trace: core/decoder.sv:591:19
										if (~CVA6Cfg[16552])
											// Trace: core/decoder.sv:592:21
											illegal_instr = 1'b1;
										(* full_case, parallel_case *)
										case (instr[13-:2])
											2'b00: begin
												// Trace: core/decoder.sv:597:23
												if (~CVA6Cfg[16437])
													// Trace: core/decoder.sv:598:25
													illegal_instr = 1'b1;
												if (instr[14])
													// Trace: core/decoder.sv:600:25
													illegal_instr = 1'b1;
											end
											2'b01:
												// Trace: core/decoder.sv:603:23
												if (~CVA6Cfg[16435])
													// Trace: core/decoder.sv:604:25
													illegal_instr = 1'b1;
											2'b10:
												// Trace: core/decoder.sv:607:23
												if (~CVA6Cfg[16436])
													// Trace: core/decoder.sv:608:25
													illegal_instr = 1'b1;
											2'b11:
												// Trace: core/decoder.sv:611:23
												if (~CVA6Cfg[16434])
													// Trace: core/decoder.sv:612:25
													illegal_instr = 1'b1;
											default:
												// Trace: core/decoder.sv:614:30
												illegal_instr = 1'b1;
										endcase
									end
									5'b11001: begin
										// Trace: core/decoder.sv:618:19
										instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd134;
										// Trace: core/decoder.sv:619:19
										imm_select = 4'd2;
										// Trace: core/decoder.sv:620:19
										if (~CVA6Cfg[16552])
											// Trace: core/decoder.sv:621:21
											illegal_instr = 1'b1;
										(* full_case, parallel_case *)
										case (instr[13-:2])
											2'b00:
												// Trace: core/decoder.sv:625:30
												illegal_instr = 1'b1;
											2'b01:
												// Trace: core/decoder.sv:626:30
												illegal_instr = 1'b1;
											2'b10:
												// Trace: core/decoder.sv:627:30
												illegal_instr = 1'b1;
											2'b11:
												// Trace: core/decoder.sv:629:23
												if (~CVA6Cfg[16434])
													// Trace: core/decoder.sv:630:25
													illegal_instr = 1'b1;
											default:
												// Trace: core/decoder.sv:632:30
												illegal_instr = 1'b1;
										endcase
									end
									5'b11010: begin
										// Trace: core/decoder.sv:636:19
										instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd135;
										// Trace: core/decoder.sv:637:19
										imm_select = 4'd2;
										// Trace: core/decoder.sv:638:19
										if (~CVA6Cfg[16551])
											// Trace: core/decoder.sv:639:21
											illegal_instr = 1'b1;
										(* full_case, parallel_case *)
										case (instr[13-:2])
											2'b00: begin
												// Trace: core/decoder.sv:644:23
												if (~CVA6Cfg[16437])
													// Trace: core/decoder.sv:645:25
													illegal_instr = 1'b1;
												if (instr[14])
													// Trace: core/decoder.sv:647:25
													illegal_instr = 1'b1;
											end
											2'b01:
												// Trace: core/decoder.sv:650:23
												if (~CVA6Cfg[16435])
													// Trace: core/decoder.sv:651:25
													illegal_instr = 1'b1;
											2'b10:
												// Trace: core/decoder.sv:654:23
												if (~CVA6Cfg[16436])
													// Trace: core/decoder.sv:655:25
													illegal_instr = 1'b1;
											2'b11:
												// Trace: core/decoder.sv:658:23
												if (~CVA6Cfg[16434])
													// Trace: core/decoder.sv:659:25
													illegal_instr = 1'b1;
											default:
												// Trace: core/decoder.sv:661:30
												illegal_instr = 1'b1;
										endcase
									end
									5'b11011: begin
										// Trace: core/decoder.sv:665:19
										instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd136;
										// Trace: core/decoder.sv:666:19
										imm_select = 4'd2;
										// Trace: core/decoder.sv:667:19
										if (~CVA6Cfg[16551])
											// Trace: core/decoder.sv:668:21
											illegal_instr = 1'b1;
										(* full_case, parallel_case *)
										case (instr[13-:2])
											2'b00:
												// Trace: core/decoder.sv:672:30
												illegal_instr = 1'b1;
											2'b01:
												// Trace: core/decoder.sv:673:30
												illegal_instr = 1'b1;
											2'b10:
												// Trace: core/decoder.sv:674:30
												illegal_instr = 1'b1;
											2'b11:
												// Trace: core/decoder.sv:676:23
												if (~CVA6Cfg[16434])
													// Trace: core/decoder.sv:677:25
													illegal_instr = 1'b1;
											default:
												// Trace: core/decoder.sv:679:30
												illegal_instr = 1'b1;
										endcase
									end
									default:
										// Trace: core/decoder.sv:682:26
										illegal_instr = 1'b1;
								endcase
								(* full_case, parallel_case *)
								case (instr[13-:2])
									2'b00:
										if (~CVA6Cfg[16437])
											// Trace: core/decoder.sv:688:47
											illegal_instr = 1'b1;
									2'b01:
										if (~CVA6Cfg[16435])
											// Trace: core/decoder.sv:689:51
											illegal_instr = 1'b1;
									2'b10:
										if (~CVA6Cfg[16436])
											// Trace: core/decoder.sv:690:48
											illegal_instr = 1'b1;
									2'b11:
										if (~CVA6Cfg[16434])
											// Trace: core/decoder.sv:691:47
											illegal_instr = 1'b1;
									default:
										// Trace: core/decoder.sv:692:26
										illegal_instr = 1'b1;
								endcase
								if (~allow_replication & instr[14])
									// Trace: core/decoder.sv:696:60
									illegal_instr = 1'b1;
								if (check_fprm) begin
									begin
										// Trace: core/decoder.sv:700:17
										(* full_case, parallel_case *)
										if ((3'b000 <= frm_i) && (3'b100 >= frm_i))
											;
										else
											// Trace: core/decoder.sv:702:28
											illegal_instr = 1'b1;
									end
								end
							end
							else
								// Trace: core/decoder.sv:707:15
								illegal_instr = 1'b1;
						end
					end
					else begin
						// Trace: core/decoder.sv:714:13
						if (CVA6Cfg[16546])
							// Trace: core/decoder.sv:715:15
							instruction_o[27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = ((instr[31-:7] == 7'b0000001) || ((instr[31-:7] == 7'b0000101) && !instr[14]) ? 4'd5 : 4'd3);
						else
							// Trace: core/decoder.sv:717:15
							instruction_o[27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = (instr[31-:7] == 7'b0000001 ? 4'd5 : 4'd3);
						// Trace: core/decoder.sv:719:13
						instruction_o[15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[19-:5];
						// Trace: core/decoder.sv:720:13
						instruction_o[10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[24-:5];
						// Trace: core/decoder.sv:721:13
						instruction_o[5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[11-:5];
						(* full_case, parallel_case *)
						case ({instr[31-:7], instr[14-:3]})
							10'b0000000000:
								// Trace: core/decoder.sv:726:39
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd0;
							10'b0100000000:
								// Trace: core/decoder.sv:727:39
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd1;
							10'b0000000010:
								// Trace: core/decoder.sv:728:39
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd21;
							10'b0000000011:
								// Trace: core/decoder.sv:732:15
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd22;
							10'b0000000100:
								// Trace: core/decoder.sv:733:39
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd4;
							10'b0000000110:
								// Trace: core/decoder.sv:734:39
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd5;
							10'b0000000111:
								// Trace: core/decoder.sv:735:39
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd6;
							10'b0000000001:
								// Trace: core/decoder.sv:736:39
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd9;
							10'b0000000101:
								// Trace: core/decoder.sv:737:39
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd8;
							10'b0100000101:
								// Trace: core/decoder.sv:738:39
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd7;
							10'b0000001000:
								// Trace: core/decoder.sv:740:39
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd83;
							10'b0000001001:
								// Trace: core/decoder.sv:741:39
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd84;
							10'b0000001010:
								// Trace: core/decoder.sv:742:39
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd86;
							10'b0000001011:
								// Trace: core/decoder.sv:743:39
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd85;
							10'b0000001100:
								// Trace: core/decoder.sv:744:39
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd88;
							10'b0000001101:
								// Trace: core/decoder.sv:745:39
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd89;
							10'b0000001110:
								// Trace: core/decoder.sv:746:39
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd92;
							10'b0000001111:
								// Trace: core/decoder.sv:747:39
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd93;
							default:
								// Trace: core/decoder.sv:749:17
								illegal_instr_non_bm = 1'b1;
						endcase
						if (CVA6Cfg[16546])
							// Trace: core/decoder.sv:753:15
							(* full_case, parallel_case *)
							case ({instr[31-:7], instr[14-:3]})
								10'b0100000111:
									// Trace: core/decoder.sv:757:41
									instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd178;
								10'b0100000110:
									// Trace: core/decoder.sv:758:41
									instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd179;
								10'b0100000100:
									// Trace: core/decoder.sv:759:41
									instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd180;
								10'b0010000010:
									// Trace: core/decoder.sv:761:41
									instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd175;
								10'b0010000100:
									// Trace: core/decoder.sv:762:41
									instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd176;
								10'b0010000110:
									// Trace: core/decoder.sv:763:41
									instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd177;
								10'b0000101110:
									// Trace: core/decoder.sv:765:41
									instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd166;
								10'b0000101111:
									// Trace: core/decoder.sv:766:41
									instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd167;
								10'b0000101100:
									// Trace: core/decoder.sv:767:41
									instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd168;
								10'b0000101101:
									// Trace: core/decoder.sv:768:41
									instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd169;
								10'b0100100001:
									// Trace: core/decoder.sv:770:41
									instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd158;
								10'b0100100101:
									// Trace: core/decoder.sv:771:41
									instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd160;
								10'b0110100001:
									// Trace: core/decoder.sv:772:41
									instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd162;
								10'b0010100001:
									// Trace: core/decoder.sv:773:41
									instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd164;
								10'b0000101001:
									// Trace: core/decoder.sv:775:41
									instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd155;
								10'b0000101011:
									// Trace: core/decoder.sv:776:41
									instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd156;
								10'b0000101010:
									// Trace: core/decoder.sv:777:41
									instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd157;
								10'b0110000001:
									// Trace: core/decoder.sv:779:41
									instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd140;
								10'b0110000101:
									// Trace: core/decoder.sv:780:41
									instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd142;
								10'b0000100100:
									// Trace: core/decoder.sv:785:19
									if (!CVA6Cfg[16973] && (instr[24:20] == 5'b00000))
										// Trace: core/decoder.sv:786:21
										instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd148;
									else
										// Trace: core/decoder.sv:787:24
										illegal_instr_bm = 1'b1;
								default:
									// Trace: core/decoder.sv:790:19
									illegal_instr_bm = 1'b1;
							endcase
						if (CVA6Cfg[16538])
							// Trace: core/decoder.sv:795:15
							(* full_case, parallel_case *)
							case ({instr[31-:7], instr[14-:3]})
								10'b0000111101:
									// Trace: core/decoder.sv:799:41
									instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd186;
								10'b0000111111:
									// Trace: core/decoder.sv:800:41
									instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd187;
								default:
									// Trace: core/decoder.sv:802:19
									illegal_instr_zic = 1'b1;
							endcase
						(* full_case, parallel_case *)
						case ({CVA6Cfg[16546], CVA6Cfg[16538]})
							2'b00:
								// Trace: core/decoder.sv:810:22
								illegal_instr = illegal_instr_non_bm;
							2'b01:
								// Trace: core/decoder.sv:811:22
								illegal_instr = illegal_instr_non_bm & illegal_instr_zic;
							2'b10:
								// Trace: core/decoder.sv:812:22
								illegal_instr = illegal_instr_non_bm & illegal_instr_bm;
							2'b11:
								// Trace: core/decoder.sv:813:22
								illegal_instr = (illegal_instr_non_bm & illegal_instr_bm) & illegal_instr_zic;
						endcase
					end
				riscv_OpcodeOp32: begin
					// Trace: core/decoder.sv:822:11
					instruction_o[27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = (instr[31-:7] == 7'b0000001 ? 4'd5 : 4'd3);
					// Trace: core/decoder.sv:823:11
					instruction_o[15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[19-:5];
					// Trace: core/decoder.sv:824:11
					instruction_o[10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[24-:5];
					// Trace: core/decoder.sv:825:11
					instruction_o[5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[11-:5];
					// Trace: core/decoder.sv:826:11
					if (CVA6Cfg[16973]) begin
						// Trace: core/decoder.sv:827:13
						(* full_case, parallel_case *)
						case ({instr[31-:7], instr[14-:3]})
							10'b0000000000:
								// Trace: core/decoder.sv:830:39
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd2;
							10'b0100000000:
								// Trace: core/decoder.sv:831:39
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd3;
							10'b0000000001:
								// Trace: core/decoder.sv:832:39
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd11;
							10'b0000000101:
								// Trace: core/decoder.sv:833:39
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd10;
							10'b0100000101:
								// Trace: core/decoder.sv:834:39
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd12;
							10'b0000001000:
								// Trace: core/decoder.sv:836:39
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd87;
							10'b0000001100:
								// Trace: core/decoder.sv:837:39
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd90;
							10'b0000001101:
								// Trace: core/decoder.sv:838:39
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd91;
							10'b0000001110:
								// Trace: core/decoder.sv:839:39
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd94;
							10'b0000001111:
								// Trace: core/decoder.sv:840:39
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd95;
							default:
								// Trace: core/decoder.sv:841:24
								illegal_instr_non_bm = 1'b1;
						endcase
						if (CVA6Cfg[16546]) begin
							// Trace: core/decoder.sv:844:15
							(* full_case, parallel_case *)
							case ({instr[31-:7], instr[14-:3]})
								10'b0010000010:
									// Trace: core/decoder.sv:848:40
									instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd170;
								10'b0010000100:
									// Trace: core/decoder.sv:849:40
									instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd171;
								10'b0010000110:
									// Trace: core/decoder.sv:850:40
									instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd172;
								10'b0000100000:
									// Trace: core/decoder.sv:852:40
									instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd173;
								10'b0110000001:
									// Trace: core/decoder.sv:854:40
									instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd141;
								10'b0110000101:
									// Trace: core/decoder.sv:855:40
									instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd145;
								10'b0000100100:
									// Trace: core/decoder.sv:859:19
									if (instr[24:20] == 5'b00000)
										// Trace: core/decoder.sv:860:21
										instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd148;
									else
										// Trace: core/decoder.sv:862:21
										illegal_instr_bm = 1'b1;
								default:
									// Trace: core/decoder.sv:864:26
									illegal_instr_bm = 1'b1;
							endcase
							// Trace: core/decoder.sv:866:15
							illegal_instr = illegal_instr_non_bm & illegal_instr_bm;
						end
						else
							// Trace: core/decoder.sv:868:15
							illegal_instr = illegal_instr_non_bm;
					end
					else
						// Trace: core/decoder.sv:870:20
						illegal_instr = 1'b1;
				end
				riscv_OpcodeOpImm: begin
					// Trace: core/decoder.sv:876:11
					instruction_o[27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 4'd3;
					// Trace: core/decoder.sv:877:11
					imm_select = 4'd1;
					// Trace: core/decoder.sv:878:11
					instruction_o[15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[19-:5];
					// Trace: core/decoder.sv:879:11
					instruction_o[5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[11-:5];
					// Trace: core/decoder.sv:880:11
					(* full_case, parallel_case *)
					case (instr[14-:3])
						3'b000:
							// Trace: core/decoder.sv:881:21
							instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd0;
						3'b010:
							// Trace: core/decoder.sv:882:21
							instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd21;
						3'b011:
							// Trace: core/decoder.sv:884:13
							instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd22;
						3'b100:
							// Trace: core/decoder.sv:885:21
							instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd4;
						3'b110:
							// Trace: core/decoder.sv:886:21
							instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd5;
						3'b111:
							// Trace: core/decoder.sv:887:21
							instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd6;
						3'b001: begin
							// Trace: core/decoder.sv:890:15
							instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd9;
							// Trace: core/decoder.sv:891:15
							if (instr[31:26] != 6'b000000)
								// Trace: core/decoder.sv:891:47
								illegal_instr_non_bm = 1'b1;
							if ((instr[25] != 1'b0) && (CVA6Cfg[17102-:32] == 32))
								// Trace: core/decoder.sv:892:66
								illegal_instr_non_bm = 1'b1;
						end
						3'b101: begin
							// Trace: core/decoder.sv:896:15
							if (instr[31:26] == 6'b000000)
								// Trace: core/decoder.sv:897:17
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd8;
							else if (instr[31:26] == 6'b010000)
								// Trace: core/decoder.sv:899:17
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd7;
							else
								// Trace: core/decoder.sv:900:20
								illegal_instr_non_bm = 1'b1;
							if ((instr[25] != 1'b0) && (CVA6Cfg[17102-:32] == 32))
								// Trace: core/decoder.sv:901:66
								illegal_instr_non_bm = 1'b1;
						end
					endcase
					if (CVA6Cfg[16546]) begin
						// Trace: core/decoder.sv:905:13
						(* full_case, parallel_case *)
						case (instr[14-:3])
							3'b001:
								// Trace: core/decoder.sv:907:17
								if (instr[31:25] == 7'b0110000) begin
									begin
										// Trace: core/decoder.sv:908:19
										if (instr[24:20] == 5'b00100)
											// Trace: core/decoder.sv:908:55
											instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd146;
										else if (instr[24:20] == 5'b00101)
											// Trace: core/decoder.sv:909:60
											instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd147;
										else if (instr[24:20] == 5'b00010)
											// Trace: core/decoder.sv:910:60
											instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd149;
										else if (instr[24:20] == 5'b00000)
											// Trace: core/decoder.sv:911:60
											instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd151;
										else if (instr[24:20] == 5'b00001)
											// Trace: core/decoder.sv:912:60
											instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd153;
										else
											// Trace: core/decoder.sv:913:24
											illegal_instr_bm = 1'b1;
									end
								end
								else if (instr[31:26] == 6'b010010)
									// Trace: core/decoder.sv:914:63
									instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd159;
								else if (instr[31:26] == 6'b011010)
									// Trace: core/decoder.sv:915:59
									instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd163;
								else if (instr[31:26] == 6'b001010)
									// Trace: core/decoder.sv:916:59
									instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd165;
								else
									// Trace: core/decoder.sv:917:22
									illegal_instr_bm = 1'b1;
							3'b101:
								// Trace: core/decoder.sv:920:17
								if (instr[31:20] == 12'b001010000111)
									// Trace: core/decoder.sv:920:61
									instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd138;
								else if (CVA6Cfg[16973] && (instr[31:20] == 12'b011010111000))
									// Trace: core/decoder.sv:922:19
									instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd139;
								else if (instr[31:20] == 12'b011010011000)
									// Trace: core/decoder.sv:924:19
									instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd139;
								else if (instr[31:26] == 6'b010010)
									// Trace: core/decoder.sv:925:60
									instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd161;
								else if (instr[31:26] == 6'b011000)
									// Trace: core/decoder.sv:926:60
									instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd143;
								else
									// Trace: core/decoder.sv:927:22
									illegal_instr_bm = 1'b1;
							default:
								// Trace: core/decoder.sv:929:24
								illegal_instr_bm = 1'b1;
						endcase
						// Trace: core/decoder.sv:931:13
						illegal_instr = illegal_instr_non_bm & illegal_instr_bm;
					end
					else
						// Trace: core/decoder.sv:933:13
						illegal_instr = illegal_instr_non_bm;
				end
				riscv_OpcodeOpImm32: begin
					// Trace: core/decoder.sv:941:11
					instruction_o[27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 4'd3;
					// Trace: core/decoder.sv:942:11
					imm_select = 4'd1;
					// Trace: core/decoder.sv:943:11
					instruction_o[15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[19-:5];
					// Trace: core/decoder.sv:944:11
					instruction_o[5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[11-:5];
					// Trace: core/decoder.sv:945:11
					if (CVA6Cfg[16973]) begin
						// Trace: core/decoder.sv:946:13
						(* full_case, parallel_case *)
						case (instr[14-:3])
							3'b000:
								// Trace: core/decoder.sv:947:24
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd2;
							3'b001: begin
								// Trace: core/decoder.sv:949:17
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd11;
								// Trace: core/decoder.sv:950:17
								if (instr[31:25] != 7'b0000000)
									// Trace: core/decoder.sv:950:49
									illegal_instr_non_bm = 1'b1;
							end
							3'b101:
								// Trace: core/decoder.sv:953:17
								if (instr[31:25] == 7'b0000000)
									// Trace: core/decoder.sv:954:19
									instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd10;
								else if (instr[31:25] == 7'b0100000)
									// Trace: core/decoder.sv:956:19
									instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd12;
								else
									// Trace: core/decoder.sv:957:22
									illegal_instr_non_bm = 1'b1;
							default:
								// Trace: core/decoder.sv:959:24
								illegal_instr_non_bm = 1'b1;
						endcase
						if (CVA6Cfg[16546]) begin
							// Trace: core/decoder.sv:962:15
							(* full_case, parallel_case *)
							case (instr[14-:3])
								3'b001:
									// Trace: core/decoder.sv:964:19
									if (instr[31:25] == 7'b0110000) begin
										begin
											// Trace: core/decoder.sv:965:21
											if (instr[21:20] == 2'b10)
												// Trace: core/decoder.sv:965:54
												instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd150;
											else if (instr[21:20] == 2'b00)
												// Trace: core/decoder.sv:966:59
												instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd152;
											else if (instr[21:20] == 2'b01)
												// Trace: core/decoder.sv:967:59
												instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd154;
											else
												// Trace: core/decoder.sv:968:26
												illegal_instr_bm = 1'b1;
										end
									end
									else if (instr[31:26] == 6'b000010)
										// Trace: core/decoder.sv:970:21
										instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd174;
									else
										// Trace: core/decoder.sv:971:28
										illegal_instr_bm = 1'b1;
								3'b101:
									// Trace: core/decoder.sv:974:19
									if (instr[31:25] == 7'b0110000)
										// Trace: core/decoder.sv:974:58
										instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd144;
									else
										// Trace: core/decoder.sv:975:24
										illegal_instr_bm = 1'b1;
								default:
									// Trace: core/decoder.sv:977:26
									illegal_instr_bm = 1'b1;
							endcase
							// Trace: core/decoder.sv:979:15
							illegal_instr = illegal_instr_non_bm & illegal_instr_bm;
						end
						else
							// Trace: core/decoder.sv:981:15
							illegal_instr = illegal_instr_non_bm;
					end
					else
						// Trace: core/decoder.sv:984:20
						illegal_instr = 1'b1;
				end
				riscv_OpcodeStore: begin
					// Trace: core/decoder.sv:990:11
					instruction_o[27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 4'd2;
					// Trace: core/decoder.sv:991:11
					imm_select = 4'd2;
					// Trace: core/decoder.sv:992:11
					instruction_o[15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[19-:5];
					// Trace: core/decoder.sv:993:11
					instruction_o[10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[24-:5];
					// Trace: core/decoder.sv:995:11
					(* full_case, parallel_case *)
					case (instr[14-:3])
						3'b000:
							// Trace: core/decoder.sv:996:21
							instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd46;
						3'b001:
							// Trace: core/decoder.sv:997:21
							instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd44;
						3'b010:
							// Trace: core/decoder.sv:998:21
							instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd41;
						3'b011:
							if (CVA6Cfg[17102-:32] == 64)
								// Trace: core/decoder.sv:1000:37
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd38;
							else
								// Trace: core/decoder.sv:1001:18
								illegal_instr = 1'b1;
						default:
							// Trace: core/decoder.sv:1002:22
							illegal_instr = 1'b1;
					endcase
					if (CVA6Cfg[16543]) begin
						// Trace: core/decoder.sv:1005:13
						tinst = {7'b0000000, instr[24-:5], 5'b00000, instr[14-:3], 5'b00000, instr[6-:7]};
						// Trace: core/decoder.sv:1006:13
						tinst[1] = (is_compressed_i ? 1'b0 : 'b1);
					end
				end
				riscv_OpcodeLoad: begin
					// Trace: core/decoder.sv:1011:11
					instruction_o[27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 4'd1;
					// Trace: core/decoder.sv:1012:11
					imm_select = 4'd1;
					// Trace: core/decoder.sv:1013:11
					instruction_o[15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[19-:5];
					// Trace: core/decoder.sv:1014:11
					instruction_o[5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[11-:5];
					// Trace: core/decoder.sv:1016:11
					(* full_case, parallel_case *)
					case (instr[14-:3])
						3'b000:
							// Trace: core/decoder.sv:1017:21
							instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd45;
						3'b001:
							// Trace: core/decoder.sv:1018:21
							instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd42;
						3'b010:
							// Trace: core/decoder.sv:1019:21
							instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd39;
						3'b100:
							// Trace: core/decoder.sv:1020:21
							instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd47;
						3'b101:
							// Trace: core/decoder.sv:1021:21
							instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd43;
						3'b110:
							if (CVA6Cfg[17102-:32] == 64)
								// Trace: core/decoder.sv:1023:37
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd40;
							else
								// Trace: core/decoder.sv:1024:18
								illegal_instr = 1'b1;
						3'b011:
							if (CVA6Cfg[17102-:32] == 64)
								// Trace: core/decoder.sv:1026:37
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd37;
							else
								// Trace: core/decoder.sv:1027:18
								illegal_instr = 1'b1;
						default:
							// Trace: core/decoder.sv:1028:22
							illegal_instr = 1'b1;
					endcase
					if (CVA6Cfg[16543]) begin
						// Trace: core/decoder.sv:1031:13
						tinst = {17'b00000000000000000, instr[14-:3], instr[11-:5], instr[6-:7]};
						// Trace: core/decoder.sv:1032:13
						tinst[1] = (is_compressed_i ? 1'b0 : 'b1);
					end
				end
				riscv_OpcodeStoreFp:
					// Trace: core/decoder.sv:1040:11
					if ((CVA6Cfg[16471] && (fs_i != 2'b00)) && ((CVA6Cfg[16543] && (!v_i || (vfs_i != 2'b00))) || !CVA6Cfg[16543])) begin
						// Trace: core/decoder.sv:1041:13
						instruction_o[27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 4'd2;
						// Trace: core/decoder.sv:1042:13
						imm_select = 4'd2;
						// Trace: core/decoder.sv:1043:13
						instruction_o[15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[19-:5];
						// Trace: core/decoder.sv:1044:13
						instruction_o[10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[24-:5];
						// Trace: core/decoder.sv:1046:13
						(* full_case, parallel_case *)
						case (instr[14-:3])
							3'b000:
								if (CVA6Cfg[16548])
									// Trace: core/decoder.sv:1049:32
									instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd103;
								else
									// Trace: core/decoder.sv:1050:20
									illegal_instr = 1'b1;
							3'b001:
								if (CVA6Cfg[16550] | CVA6Cfg[16549])
									// Trace: core/decoder.sv:1052:51
									instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd102;
								else
									// Trace: core/decoder.sv:1053:20
									illegal_instr = 1'b1;
							3'b010:
								if (CVA6Cfg[16552])
									// Trace: core/decoder.sv:1055:32
									instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd101;
								else
									// Trace: core/decoder.sv:1056:20
									illegal_instr = 1'b1;
							3'b011:
								if (CVA6Cfg[16551])
									// Trace: core/decoder.sv:1058:32
									instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd100;
								else
									// Trace: core/decoder.sv:1059:20
									illegal_instr = 1'b1;
							default:
								// Trace: core/decoder.sv:1060:24
								illegal_instr = 1'b1;
						endcase
						if (CVA6Cfg[16543]) begin
							// Trace: core/decoder.sv:1063:15
							tinst = {7'b0000000, instr[24-:5], 5'b00000, instr[14-:3], 5'b00000, instr[6-:7]};
							// Trace: core/decoder.sv:1064:15
							tinst[1] = (is_compressed_i ? 1'b0 : 'b1);
						end
					end
					else
						// Trace: core/decoder.sv:1066:20
						illegal_instr = 1'b1;
				riscv_OpcodeLoadFp:
					// Trace: core/decoder.sv:1070:11
					if ((CVA6Cfg[16471] && (fs_i != 2'b00)) && ((CVA6Cfg[16543] && (!v_i || (vfs_i != 2'b00))) || !CVA6Cfg[16543])) begin
						// Trace: core/decoder.sv:1071:13
						instruction_o[27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 4'd1;
						// Trace: core/decoder.sv:1072:13
						imm_select = 4'd1;
						// Trace: core/decoder.sv:1073:13
						instruction_o[15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[19-:5];
						// Trace: core/decoder.sv:1074:13
						instruction_o[5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[11-:5];
						// Trace: core/decoder.sv:1076:13
						(* full_case, parallel_case *)
						case (instr[14-:3])
							3'b000:
								if (CVA6Cfg[16548])
									// Trace: core/decoder.sv:1079:32
									instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd99;
								else
									// Trace: core/decoder.sv:1080:20
									illegal_instr = 1'b1;
							3'b001:
								if (CVA6Cfg[16550] | CVA6Cfg[16549])
									// Trace: core/decoder.sv:1082:51
									instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd98;
								else
									// Trace: core/decoder.sv:1083:20
									illegal_instr = 1'b1;
							3'b010:
								if (CVA6Cfg[16552])
									// Trace: core/decoder.sv:1085:32
									instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd97;
								else
									// Trace: core/decoder.sv:1086:20
									illegal_instr = 1'b1;
							3'b011:
								if (CVA6Cfg[16551])
									// Trace: core/decoder.sv:1088:32
									instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd96;
								else
									// Trace: core/decoder.sv:1089:20
									illegal_instr = 1'b1;
							default:
								// Trace: core/decoder.sv:1090:24
								illegal_instr = 1'b1;
						endcase
						if (CVA6Cfg[16543]) begin
							// Trace: core/decoder.sv:1093:15
							tinst = {17'b00000000000000000, instr[14-:3], instr[11-:5], instr[6-:7]};
							// Trace: core/decoder.sv:1094:15
							tinst[1] = (is_compressed_i ? 1'b0 : 'b1);
						end
					end
					else
						// Trace: core/decoder.sv:1096:20
						illegal_instr = 1'b1;
				riscv_OpcodeMadd, riscv_OpcodeMsub, riscv_OpcodeNmsub, riscv_OpcodeNmadd:
					// Trace: core/decoder.sv:1103:11
					if ((CVA6Cfg[16471] && (fs_i != 2'b00)) && ((CVA6Cfg[16543] && (!v_i || (vfs_i != 2'b00))) || !CVA6Cfg[16543])) begin
						// Trace: core/decoder.sv:1104:13
						instruction_o[27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 4'd7;
						// Trace: core/decoder.sv:1105:13
						instruction_o[15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[19-:5];
						// Trace: core/decoder.sv:1106:13
						instruction_o[10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[24-:5];
						// Trace: core/decoder.sv:1107:13
						instruction_o[5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[11-:5];
						// Trace: core/decoder.sv:1108:13
						imm_select = 4'd6;
						// Trace: core/decoder.sv:1109:13
						check_fprm = 1'b1;
						// Trace: core/decoder.sv:1111:13
						(* full_case, parallel_case *)
						case (instr[6-:7])
							default:
								// Trace: core/decoder.sv:1112:24
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd110;
							riscv_OpcodeMsub:
								// Trace: core/decoder.sv:1114:15
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd111;
							riscv_OpcodeNmsub:
								// Trace: core/decoder.sv:1116:15
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd112;
							riscv_OpcodeNmadd:
								// Trace: core/decoder.sv:1118:15
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd113;
						endcase
						(* full_case, parallel_case *)
						case (instr[26-:2])
							2'b00:
								if (~CVA6Cfg[16552])
									// Trace: core/decoder.sv:1124:42
									illegal_instr = 1'b1;
							2'b01:
								if (~CVA6Cfg[16551])
									// Trace: core/decoder.sv:1125:42
									illegal_instr = 1'b1;
							2'b10:
								if (~CVA6Cfg[16550] & ~CVA6Cfg[16549])
									// Trace: core/decoder.sv:1126:62
									illegal_instr = 1'b1;
							2'b11:
								if (~CVA6Cfg[16548])
									// Trace: core/decoder.sv:1127:42
									illegal_instr = 1'b1;
							default:
								// Trace: core/decoder.sv:1128:24
								illegal_instr = 1'b1;
						endcase
						if (check_fprm) begin
							begin
								// Trace: core/decoder.sv:1133:15
								(* full_case, parallel_case *)
								if ((3'b000 <= instr[14-:3]) && (3'b100 >= instr[14-:3]))
									;
								else if (instr[14-:3] == 3'b101) begin
									// Trace: core/decoder.sv:1136:19
									if (~CVA6Cfg[16549] || (instr[26-:2] != 2'b10))
										// Trace: core/decoder.sv:1136:70
										illegal_instr = 1'b1;
									(* full_case, parallel_case *)
									if ((3'b000 <= frm_i) && (3'b100 >= frm_i))
										;
									else
										// Trace: core/decoder.sv:1139:30
										illegal_instr = 1'b1;
								end
								else if (instr[14-:3] == 3'b111) begin
									begin
										// Trace: core/decoder.sv:1144:19
										(* full_case, parallel_case *)
										if ((3'b000 <= frm_i) && (3'b100 >= frm_i))
											;
										else
											// Trace: core/decoder.sv:1146:30
											illegal_instr = 1'b1;
									end
								end
								else
									// Trace: core/decoder.sv:1149:36
									illegal_instr = 1'b1;
							end
						end
					end
					else
						// Trace: core/decoder.sv:1153:13
						illegal_instr = 1'b1;
				riscv_OpcodeOpFp:
					// Trace: core/decoder.sv:1158:11
					if ((CVA6Cfg[16471] && (fs_i != 2'b00)) && ((CVA6Cfg[16543] && (!v_i || (vfs_i != 2'b00))) || !CVA6Cfg[16543])) begin
						// Trace: core/decoder.sv:1159:13
						instruction_o[27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 4'd7;
						// Trace: core/decoder.sv:1160:13
						instruction_o[15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[19-:5];
						// Trace: core/decoder.sv:1161:13
						instruction_o[10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[24-:5];
						// Trace: core/decoder.sv:1162:13
						instruction_o[5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[11-:5];
						// Trace: core/decoder.sv:1163:13
						check_fprm = 1'b1;
						// Trace: core/decoder.sv:1165:13
						(* full_case, parallel_case *)
						case (instr[31-:5])
							5'b00000: begin
								// Trace: core/decoder.sv:1167:17
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd104;
								// Trace: core/decoder.sv:1168:17
								instruction_o[15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 1'sb0;
								// Trace: core/decoder.sv:1169:17
								instruction_o[10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[19-:5];
								// Trace: core/decoder.sv:1170:17
								imm_select = 4'd1;
							end
							5'b00001: begin
								// Trace: core/decoder.sv:1173:17
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd105;
								// Trace: core/decoder.sv:1174:17
								instruction_o[15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 1'sb0;
								// Trace: core/decoder.sv:1175:17
								instruction_o[10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[19-:5];
								// Trace: core/decoder.sv:1176:17
								imm_select = 4'd1;
							end
							5'b00010:
								// Trace: core/decoder.sv:1178:25
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd106;
							5'b00011:
								// Trace: core/decoder.sv:1179:25
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd107;
							5'b01011: begin
								// Trace: core/decoder.sv:1181:17
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd109;
								// Trace: core/decoder.sv:1183:17
								if (instr[24-:5] != 5'b00000)
									// Trace: core/decoder.sv:1183:51
									illegal_instr = 1'b1;
							end
							5'b00100: begin
								// Trace: core/decoder.sv:1186:17
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd117;
								// Trace: core/decoder.sv:1187:17
								check_fprm = 1'b0;
								// Trace: core/decoder.sv:1188:17
								if (CVA6Cfg[16549]) begin
									begin
										// Trace: core/decoder.sv:1189:19
										if (!(|{(3'b000 <= instr[14-:3]) && (3'b010 >= instr[14-:3]), (3'b100 <= instr[14-:3]) && (3'b110 >= instr[14-:3])}))
											// Trace: core/decoder.sv:1190:21
											illegal_instr = 1'b1;
									end
								end
								else
									// Trace: core/decoder.sv:1192:19
									if (!((3'b000 <= instr[14-:3]) && (3'b010 >= instr[14-:3])))
										// Trace: core/decoder.sv:1192:70
										illegal_instr = 1'b1;
							end
							5'b00101: begin
								// Trace: core/decoder.sv:1196:17
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd108;
								// Trace: core/decoder.sv:1197:17
								check_fprm = 1'b0;
								// Trace: core/decoder.sv:1198:17
								if (CVA6Cfg[16549]) begin
									begin
										// Trace: core/decoder.sv:1199:19
										if (!(|{(3'b000 <= instr[14-:3]) && (3'b001 >= instr[14-:3]), (3'b100 <= instr[14-:3]) && (3'b101 >= instr[14-:3])}))
											// Trace: core/decoder.sv:1200:21
											illegal_instr = 1'b1;
									end
								end
								else
									// Trace: core/decoder.sv:1202:19
									if (!((3'b000 <= instr[14-:3]) && (3'b001 >= instr[14-:3])))
										// Trace: core/decoder.sv:1202:70
										illegal_instr = 1'b1;
							end
							5'b01000: begin
								// Trace: core/decoder.sv:1206:17
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd116;
								// Trace: core/decoder.sv:1207:17
								instruction_o[10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[19-:5];
								// Trace: core/decoder.sv:1208:17
								imm_select = 4'd1;
								// Trace: core/decoder.sv:1209:17
								if (|instr[24:23])
									// Trace: core/decoder.sv:1210:19
									illegal_instr = 1'b1;
								(* full_case, parallel_case *)
								case (instr[22:20])
									3'b000:
										if (~CVA6Cfg[16552])
											// Trace: core/decoder.sv:1214:46
											illegal_instr = 1'b1;
									3'b001:
										if (~CVA6Cfg[16551])
											// Trace: core/decoder.sv:1215:46
											illegal_instr = 1'b1;
									3'b010:
										if (~CVA6Cfg[16550])
											// Trace: core/decoder.sv:1216:47
											illegal_instr = 1'b1;
									3'b110:
										if (~CVA6Cfg[16549])
											// Trace: core/decoder.sv:1217:50
											illegal_instr = 1'b1;
									3'b011:
										if (~CVA6Cfg[16548])
											// Trace: core/decoder.sv:1218:46
											illegal_instr = 1'b1;
									default:
										// Trace: core/decoder.sv:1219:28
										illegal_instr = 1'b1;
								endcase
							end
							5'b10100: begin
								// Trace: core/decoder.sv:1223:17
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd120;
								// Trace: core/decoder.sv:1224:17
								check_fprm = 1'b0;
								// Trace: core/decoder.sv:1225:17
								if (CVA6Cfg[16549]) begin
									begin
										// Trace: core/decoder.sv:1226:19
										if (!(|{(3'b000 <= instr[14-:3]) && (3'b010 >= instr[14-:3]), (3'b100 <= instr[14-:3]) && (3'b110 >= instr[14-:3])}))
											// Trace: core/decoder.sv:1227:21
											illegal_instr = 1'b1;
									end
								end
								else
									// Trace: core/decoder.sv:1229:19
									if (!((3'b000 <= instr[14-:3]) && (3'b010 >= instr[14-:3])))
										// Trace: core/decoder.sv:1229:70
										illegal_instr = 1'b1;
							end
							5'b11000: begin
								// Trace: core/decoder.sv:1233:17
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd114;
								// Trace: core/decoder.sv:1234:17
								imm_select = 4'd1;
								// Trace: core/decoder.sv:1235:17
								if (|instr[24:22])
									// Trace: core/decoder.sv:1236:19
									illegal_instr = 1'b1;
							end
							5'b11010: begin
								// Trace: core/decoder.sv:1239:17
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd115;
								// Trace: core/decoder.sv:1240:17
								imm_select = 4'd1;
								// Trace: core/decoder.sv:1241:17
								if (|instr[24:22])
									// Trace: core/decoder.sv:1242:19
									illegal_instr = 1'b1;
							end
							5'b11100: begin
								// Trace: core/decoder.sv:1245:17
								instruction_o[10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[19-:5];
								// Trace: core/decoder.sv:1246:17
								check_fprm = 1'b0;
								// Trace: core/decoder.sv:1247:17
								if ((instr[14-:3] == 3'b000) || (CVA6Cfg[16549] && (instr[14-:3] == 3'b100)))
									// Trace: core/decoder.sv:1248:19
									instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd118;
								else if ((instr[14-:3] == 3'b001) || (CVA6Cfg[16549] && (instr[14-:3] == 3'b101)))
									// Trace: core/decoder.sv:1250:19
									instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd121;
								else
									// Trace: core/decoder.sv:1251:22
									illegal_instr = 1'b1;
								if (instr[24-:5] != 5'b00000)
									// Trace: core/decoder.sv:1253:51
									illegal_instr = 1'b1;
							end
							5'b11110: begin
								// Trace: core/decoder.sv:1256:17
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd119;
								// Trace: core/decoder.sv:1257:17
								instruction_o[10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[19-:5];
								// Trace: core/decoder.sv:1258:17
								check_fprm = 1'b0;
								// Trace: core/decoder.sv:1259:17
								if (!((instr[14-:3] == 3'b000) || (CVA6Cfg[16549] && (instr[14-:3] == 3'b100))))
									// Trace: core/decoder.sv:1260:19
									illegal_instr = 1'b1;
								if (instr[24-:5] != 5'b00000)
									// Trace: core/decoder.sv:1262:51
									illegal_instr = 1'b1;
							end
							default:
								// Trace: core/decoder.sv:1264:25
								illegal_instr = 1'b1;
						endcase
						(* full_case, parallel_case *)
						case (instr[26-:2])
							2'b00:
								if (~CVA6Cfg[16552])
									// Trace: core/decoder.sv:1270:42
									illegal_instr = 1'b1;
							2'b01:
								if (~CVA6Cfg[16551])
									// Trace: core/decoder.sv:1271:42
									illegal_instr = 1'b1;
							2'b10:
								if (~CVA6Cfg[16550] & ~CVA6Cfg[16549])
									// Trace: core/decoder.sv:1272:62
									illegal_instr = 1'b1;
							2'b11:
								if (~CVA6Cfg[16548])
									// Trace: core/decoder.sv:1273:42
									illegal_instr = 1'b1;
							default:
								// Trace: core/decoder.sv:1274:24
								illegal_instr = 1'b1;
						endcase
						if (check_fprm) begin
							begin
								// Trace: core/decoder.sv:1279:15
								(* full_case, parallel_case *)
								if ((3'b000 <= instr[14-:3]) && (3'b100 >= instr[14-:3]))
									;
								else if (instr[14-:3] == 3'b101) begin
									// Trace: core/decoder.sv:1282:19
									if (~CVA6Cfg[16549] || (instr[26-:2] != 2'b10))
										// Trace: core/decoder.sv:1282:70
										illegal_instr = 1'b1;
									(* full_case, parallel_case *)
									if ((3'b000 <= frm_i) && (3'b100 >= frm_i))
										;
									else
										// Trace: core/decoder.sv:1285:30
										illegal_instr = 1'b1;
								end
								else if (instr[14-:3] == 3'b111) begin
									begin
										// Trace: core/decoder.sv:1290:19
										(* full_case, parallel_case *)
										if ((3'b000 <= frm_i) && (3'b100 >= frm_i))
											;
										else
											// Trace: core/decoder.sv:1292:30
											illegal_instr = 1'b1;
									end
								end
								else
									// Trace: core/decoder.sv:1295:36
									illegal_instr = 1'b1;
							end
						end
					end
					else
						// Trace: core/decoder.sv:1299:13
						illegal_instr = 1'b1;
				riscv_OpcodeAmo: begin
					// Trace: core/decoder.sv:1308:11
					instruction_o[27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 4'd2;
					// Trace: core/decoder.sv:1309:11
					instruction_o[15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[19-:5];
					// Trace: core/decoder.sv:1310:11
					instruction_o[10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[24-:5];
					// Trace: core/decoder.sv:1311:11
					instruction_o[5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[11-:5];
					// Trace: core/decoder.sv:1314:11
					if (CVA6Cfg[16547] && (instr[14-:3] == 3'h2))
						// Trace: core/decoder.sv:1315:13
						(* full_case, parallel_case *)
						case (instr[31:27])
							5'h00:
								// Trace: core/decoder.sv:1316:21
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd66;
							5'h01:
								// Trace: core/decoder.sv:1317:21
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd65;
							5'h02: begin
								// Trace: core/decoder.sv:1319:17
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd61;
								// Trace: core/decoder.sv:1320:17
								if (instr[24-:5] != 0)
									// Trace: core/decoder.sv:1320:43
									illegal_instr = 1'b1;
							end
							5'h03:
								// Trace: core/decoder.sv:1322:21
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd63;
							5'h04:
								// Trace: core/decoder.sv:1323:21
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd69;
							5'h08:
								// Trace: core/decoder.sv:1324:21
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd68;
							5'h0c:
								// Trace: core/decoder.sv:1325:21
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd67;
							5'h10:
								// Trace: core/decoder.sv:1326:22
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd72;
							5'h14:
								// Trace: core/decoder.sv:1327:22
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd70;
							5'h18:
								// Trace: core/decoder.sv:1328:22
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd73;
							5'h1c:
								// Trace: core/decoder.sv:1329:22
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd71;
							default:
								// Trace: core/decoder.sv:1330:24
								illegal_instr = 1'b1;
						endcase
					else if ((CVA6Cfg[16973] && CVA6Cfg[16547]) && (instr[14-:3] == 3'h3))
						// Trace: core/decoder.sv:1334:13
						(* full_case, parallel_case *)
						case (instr[31:27])
							5'h00:
								// Trace: core/decoder.sv:1335:21
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd75;
							5'h01:
								// Trace: core/decoder.sv:1336:21
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd74;
							5'h02: begin
								// Trace: core/decoder.sv:1338:17
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd62;
								// Trace: core/decoder.sv:1339:17
								if (instr[24-:5] != 0)
									// Trace: core/decoder.sv:1339:43
									illegal_instr = 1'b1;
							end
							5'h03:
								// Trace: core/decoder.sv:1341:21
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd64;
							5'h04:
								// Trace: core/decoder.sv:1342:21
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd78;
							5'h08:
								// Trace: core/decoder.sv:1343:21
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd77;
							5'h0c:
								// Trace: core/decoder.sv:1344:21
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd76;
							5'h10:
								// Trace: core/decoder.sv:1345:22
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd81;
							5'h14:
								// Trace: core/decoder.sv:1346:22
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd79;
							5'h18:
								// Trace: core/decoder.sv:1347:22
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd82;
							5'h1c:
								// Trace: core/decoder.sv:1348:22
								instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd80;
							default:
								// Trace: core/decoder.sv:1349:24
								illegal_instr = 1'b1;
						endcase
					else
						// Trace: core/decoder.sv:1352:13
						illegal_instr = 1'b1;
					// Trace: core/decoder.sv:1354:11
					tinst = {instr[31-:5], instr[26], instr[25], instr[24-:5], 5'b00000, instr[14-:3], instr[11-:5], instr[6-:7]};
				end
				riscv_OpcodeBranch: begin
					// Trace: core/decoder.sv:1370:11
					imm_select = 4'd3;
					// Trace: core/decoder.sv:1371:11
					instruction_o[27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 4'd4;
					// Trace: core/decoder.sv:1372:11
					instruction_o[15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[19-:5];
					// Trace: core/decoder.sv:1373:11
					instruction_o[10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[24-:5];
					// Trace: core/decoder.sv:1375:11
					is_control_flow_instr_o = 1'b1;
					// Trace: core/decoder.sv:1377:11
					case (instr[14-:3])
						3'b000:
							// Trace: core/decoder.sv:1378:21
							instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd17;
						3'b001:
							// Trace: core/decoder.sv:1379:21
							instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd18;
						3'b100:
							// Trace: core/decoder.sv:1380:21
							instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd13;
						3'b101:
							// Trace: core/decoder.sv:1381:21
							instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd15;
						3'b110:
							// Trace: core/decoder.sv:1382:21
							instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd14;
						3'b111:
							// Trace: core/decoder.sv:1383:21
							instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd16;
						default: begin
							// Trace: core/decoder.sv:1385:15
							is_control_flow_instr_o = 1'b0;
							// Trace: core/decoder.sv:1386:15
							illegal_instr = 1'b1;
						end
					endcase
				end
				riscv_OpcodeJalr: begin
					// Trace: core/decoder.sv:1392:11
					instruction_o[27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 4'd4;
					// Trace: core/decoder.sv:1393:11
					instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd19;
					// Trace: core/decoder.sv:1394:11
					instruction_o[15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[19-:5];
					// Trace: core/decoder.sv:1395:11
					imm_select = 4'd1;
					// Trace: core/decoder.sv:1396:11
					instruction_o[5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[11-:5];
					// Trace: core/decoder.sv:1397:11
					is_control_flow_instr_o = 1'b1;
					// Trace: core/decoder.sv:1399:11
					if (instr[14-:3] != 3'b000)
						// Trace: core/decoder.sv:1399:43
						illegal_instr = 1'b1;
				end
				riscv_OpcodeJal: begin
					// Trace: core/decoder.sv:1403:11
					instruction_o[27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 4'd4;
					// Trace: core/decoder.sv:1404:11
					imm_select = 4'd5;
					// Trace: core/decoder.sv:1405:11
					instruction_o[5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[11-:5];
					// Trace: core/decoder.sv:1406:11
					is_control_flow_instr_o = 1'b1;
				end
				riscv_OpcodeAuipc: begin
					// Trace: core/decoder.sv:1410:11
					instruction_o[27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 4'd3;
					// Trace: core/decoder.sv:1411:11
					imm_select = 4'd4;
					// Trace: core/decoder.sv:1412:11
					instruction_o[1 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))] = 1'b1;
					// Trace: core/decoder.sv:1413:11
					instruction_o[5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[11-:5];
				end
				riscv_OpcodeLui: begin
					// Trace: core/decoder.sv:1417:11
					imm_select = 4'd4;
					// Trace: core/decoder.sv:1418:11
					instruction_o[27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 4'd3;
					// Trace: core/decoder.sv:1419:11
					instruction_o[5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[11-:5];
				end
				default:
					// Trace: core/decoder.sv:1422:18
					illegal_instr = 1'b1;
			endcase
		if (CVA6Cfg[16539]) begin
			begin
				// Trace: core/decoder.sv:1426:7
				if (~ex_i[0] && (is_illegal_i || illegal_instr)) begin
					// Trace: core/decoder.sv:1427:9
					instruction_o[27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 4'd9;
					// Trace: core/decoder.sv:1428:9
					instruction_o[15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[19-:5];
					// Trace: core/decoder.sv:1429:9
					instruction_o[10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[24-:5];
					// Trace: core/decoder.sv:1430:9
					instruction_o[5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))):(5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4] = instr[11-:5];
					// Trace: core/decoder.sv:1431:9
					instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 8'd137;
					// Trace: core/decoder.sv:1432:9
					imm_select = ((((instr[6-:7] == riscv_OpcodeMadd) || (instr[6-:7] == riscv_OpcodeMsub)) || (instr[6-:7] == riscv_OpcodeNmadd)) || (instr[6-:7] == riscv_OpcodeNmsub) ? 4'd6 : 4'd7);
				end
			end
		end
		if (CVA6Cfg[16369]) begin
			begin
				// Trace: core/decoder.sv:1442:7
				if (is_accel) begin
					// Trace: core/decoder.sv:1443:9
					instruction_o[27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = acc_instruction[27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)];
					// Trace: core/decoder.sv:1444:9
					instruction_o[0] = acc_instruction[0];
					// Trace: core/decoder.sv:1445:9
					instruction_o[15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = acc_instruction[15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)];
					// Trace: core/decoder.sv:1446:9
					instruction_o[10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = acc_instruction[10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)];
					// Trace: core/decoder.sv:1447:9
					instruction_o[5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = acc_instruction[5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)];
					// Trace: core/decoder.sv:1448:9
					instruction_o[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = acc_instruction[23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)];
					// Trace: core/decoder.sv:1449:9
					illegal_instr = acc_illegal_instr;
					// Trace: core/decoder.sv:1450:9
					is_control_flow_instr_o = acc_is_control_flow_instr;
				end
			end
		end
	end
	// Trace: core/decoder.sv:1458:3
	always @(*) begin : sign_extend
		if (_sv2v_0)
			;
		// Trace: core/decoder.sv:1459:5
		imm_i_type = {{CVA6Cfg[17102-:32] - 12 {instruction_i[31]}}, instruction_i[31:20]};
		// Trace: core/decoder.sv:1460:5
		imm_s_type = {{CVA6Cfg[17102-:32] - 12 {instruction_i[31]}}, instruction_i[31:25], instruction_i[11:7]};
		// Trace: core/decoder.sv:1463:5
		imm_sb_type = {{CVA6Cfg[17102-:32] - 13 {instruction_i[31]}}, instruction_i[31], instruction_i[7], instruction_i[30:25], instruction_i[11:8], 1'b0};
		// Trace: core/decoder.sv:1471:5
		imm_u_type = {{CVA6Cfg[17102-:32] - 32 {instruction_i[31]}}, instruction_i[31:12], 12'b000000000000};
		// Trace: core/decoder.sv:1474:5
		imm_uj_type = {{CVA6Cfg[17102-:32] - 20 {instruction_i[31]}}, instruction_i[19:12], instruction_i[20], instruction_i[30:21], 1'b0};
		// Trace: core/decoder.sv:1481:5
		imm_bi_type = {{CVA6Cfg[17102-:32] - 5 {instruction_i[24]}}, instruction_i[24:20]};
		// Trace: core/decoder.sv:1485:5
		case (imm_select)
			4'd1: begin
				// Trace: core/decoder.sv:1487:9
				instruction_o[scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))-:((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) >= (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) + 1 : ((4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + 1)] = imm_i_type;
				// Trace: core/decoder.sv:1488:9
				instruction_o[3 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))] = 1'b1;
			end
			4'd2: begin
				// Trace: core/decoder.sv:1491:9
				instruction_o[scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))-:((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) >= (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) + 1 : ((4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + 1)] = imm_s_type;
				// Trace: core/decoder.sv:1492:9
				instruction_o[3 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))] = 1'b1;
			end
			4'd3: begin
				// Trace: core/decoder.sv:1495:9
				instruction_o[scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))-:((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) >= (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) + 1 : ((4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + 1)] = imm_sb_type;
				// Trace: core/decoder.sv:1496:9
				instruction_o[3 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))] = 1'b1;
			end
			4'd4: begin
				// Trace: core/decoder.sv:1499:9
				instruction_o[scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))-:((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) >= (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) + 1 : ((4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + 1)] = imm_u_type;
				// Trace: core/decoder.sv:1500:9
				instruction_o[3 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))] = 1'b1;
			end
			4'd5: begin
				// Trace: core/decoder.sv:1503:9
				instruction_o[scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))-:((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) >= (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) + 1 : ((4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + 1)] = imm_uj_type;
				// Trace: core/decoder.sv:1504:9
				instruction_o[3 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))] = 1'b1;
			end
			4'd6: begin
				// Trace: core/decoder.sv:1508:9
				instruction_o[scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))-:((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) >= (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) + 1 : ((4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + 1)] = {{CVA6Cfg[17102-:32] - 5 {1'b0}}, instr[31-:5]};
				// Trace: core/decoder.sv:1509:9
				instruction_o[3 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))] = 1'b0;
			end
			4'd7: begin
				// Trace: core/decoder.sv:1513:9
				instruction_o[scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))-:((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) >= (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) + 1 : ((4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + 1)] = {{CVA6Cfg[17102-:32] - 5 {1'b0}}, instr[11-:5]};
				// Trace: core/decoder.sv:1514:9
				instruction_o[3 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))] = 1'b0;
			end
			default: begin
				// Trace: core/decoder.sv:1517:9
				instruction_o[scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))-:((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) >= (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) + 1 : ((4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + 1)] = {CVA6Cfg[17102-:32] {1'b0}};
				// Trace: core/decoder.sv:1518:9
				instruction_o[3 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))] = 1'b0;
			end
		endcase
		if (CVA6Cfg[16369]) begin
			begin
				// Trace: core/decoder.sv:1523:7
				if (is_accel) begin
					// Trace: core/decoder.sv:1524:9
					instruction_o[scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))-:((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) >= (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) + 1 : ((4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + 1)] = acc_instruction[scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))-:((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) >= (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) + 1 : ((4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + 1)];
					// Trace: core/decoder.sv:1525:9
					instruction_o[3 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))] = acc_instruction[3 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))];
				end
			end
		end
	end
	// Trace: core/decoder.sv:1533:3
	reg [CVA6Cfg[17102-:32] - 1:0] interrupt_cause;
	// Trace: core/decoder.sv:1536:3
	wire [1:1] sv2v_tmp_C3394;
	assign sv2v_tmp_C3394 = instruction_o[((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) : (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)];
	always @(*) instruction_o[4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))] = sv2v_tmp_C3394;
	// Trace: core/decoder.sv:1538:3
	localparam ariane_pkg_SupervisorIrq = 1;
	localparam cva6_config_pkg_CVA6ConfigXlen = 64;
	localparam riscv_XLEN = cva6_config_pkg_CVA6ConfigXlen;
	localparam [63:0] riscv_BREAKPOINT = 3;
	localparam [63:0] riscv_DEBUG_REQUEST = 24;
	localparam [63:0] riscv_ENV_CALL_MMODE = 11;
	localparam [63:0] riscv_ENV_CALL_SMODE = 9;
	localparam [63:0] riscv_ENV_CALL_UMODE = 8;
	localparam [63:0] riscv_ENV_CALL_VSMODE = 10;
	localparam [63:0] riscv_ILLEGAL_INSTR = 2;
	localparam [31:0] riscv_IRQ_HS_EXT = 12;
	localparam [31:0] riscv_IRQ_M_EXT = 11;
	localparam [31:0] riscv_IRQ_M_SOFT = 3;
	localparam [31:0] riscv_IRQ_M_TIMER = 7;
	localparam [31:0] riscv_IRQ_S_EXT = 9;
	localparam [31:0] riscv_IRQ_S_SOFT = 1;
	localparam [31:0] riscv_IRQ_S_TIMER = 5;
	localparam [31:0] riscv_IRQ_VS_EXT = 10;
	localparam [31:0] riscv_IRQ_VS_SOFT = 2;
	localparam [31:0] riscv_IRQ_VS_TIMER = 6;
	localparam [63:0] riscv_VIRTUAL_INSTRUCTION = 22;
	always @(*) begin : exception_handling
		if (_sv2v_0)
			;
		// Trace: core/decoder.sv:1539:5
		interrupt_cause = 1'sb0;
		// Trace: core/decoder.sv:1540:5
		instruction_o[((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)-:((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) >= ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5) ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) - ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)) + 1 : (((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5) - (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))) + 1)] = ex_i;
		// Trace: core/decoder.sv:1541:5
		orig_instr_o = 1'sb0;
		// Trace: core/decoder.sv:1544:5
		if (~ex_i[0]) begin
			// Trace: core/decoder.sv:1547:7
			if (CVA6Cfg[16539] || CVA6Cfg[16552])
				// Trace: core/decoder.sv:1548:9
				orig_instr_o = (is_compressed_i ? {{CVA6Cfg[17102-:32] - 16 {1'b0}}, compressed_instr_i} : {{CVA6Cfg[17102-:32] - 32 {1'b0}}, instruction_i});
			if (CVA6Cfg[15915])
				// Trace: core/decoder.sv:1550:9
				instruction_o[((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) - ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) : ((((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) + ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) + 1)) - 1)-:((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) + 1)] = (is_compressed_i ? {{CVA6Cfg[17102-:32] - 16 {1'b0}}, compressed_instr_i} : {{CVA6Cfg[17102-:32] - 32 {1'b0}}, instruction_i});
			else
				// Trace: core/decoder.sv:1551:12
				instruction_o[((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) - ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) : ((((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) + ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) + 1)) - 1)-:((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) + 1)] = 1'sb0;
			if (CVA6Cfg[16543])
				// Trace: core/decoder.sv:1552:24
				instruction_o[((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 0) : (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 3)-:32] = tinst;
			else
				// Trace: core/decoder.sv:1553:12
				instruction_o[((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 0) : (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 3)-:32] = 1'sb0;
			if (illegal_instr || is_illegal_i) begin
				// Trace: core/decoder.sv:1559:9
				if (!CVA6Cfg[16539])
					// Trace: core/decoder.sv:1559:31
					instruction_o[((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) : (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)] = 1'b1;
				// Trace: core/decoder.sv:1561:9
				instruction_o[((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) - ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) : ((((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) + ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) + 1)) - 1)-:((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) + 1)] = riscv_ILLEGAL_INSTR;
			end
			else if (CVA6Cfg[16543] && virtual_illegal_instr) begin
				// Trace: core/decoder.sv:1563:9
				instruction_o[((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) : (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)] = 1'b1;
				// Trace: core/decoder.sv:1565:9
				instruction_o[((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) - ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) : ((((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) + ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) + 1)) - 1)-:((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) + 1)] = riscv_VIRTUAL_INSTRUCTION;
			end
			else if (ecall) begin
				// Trace: core/decoder.sv:1569:9
				instruction_o[((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) : (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)] = 1'b1;
				// Trace: core/decoder.sv:1571:9
				if ((priv_lvl_i == 2'b01) && CVA6Cfg[16366])
					// Trace: core/decoder.sv:1572:11
					instruction_o[((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) - ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) : ((((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) + ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) + 1)) - 1)-:((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) + 1)] = (CVA6Cfg[16543] && v_i ? riscv_ENV_CALL_VSMODE : riscv_ENV_CALL_SMODE);
				else if ((priv_lvl_i == 2'b00) && CVA6Cfg[16365])
					// Trace: core/decoder.sv:1574:11
					instruction_o[((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) - ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) : ((((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) + ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) + 1)) - 1)-:((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) + 1)] = riscv_ENV_CALL_UMODE;
				else if (priv_lvl_i == 2'b11)
					// Trace: core/decoder.sv:1576:11
					instruction_o[((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) - ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) : ((((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) + ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) + 1)) - 1)-:((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) + 1)] = riscv_ENV_CALL_MMODE;
			end
			else if (ebreak) begin
				// Trace: core/decoder.sv:1580:9
				instruction_o[((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) : (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)] = 1'b1;
				// Trace: core/decoder.sv:1582:9
				instruction_o[((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) - ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) : ((((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) + ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) + 1)) - 1)-:((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) + 1)] = riscv_BREAKPOINT;
				// Trace: core/decoder.sv:1584:9
				if (CVA6Cfg[16543])
					// Trace: core/decoder.sv:1584:26
					instruction_o[((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 32) : (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)] = v_i;
				else
					// Trace: core/decoder.sv:1585:14
					instruction_o[((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 32) : (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)] = 1'b0;
			end
			if (CVA6Cfg[16543]) begin
				// Trace: core/decoder.sv:1596:9
				if (irq_ctrl_i[(irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + (irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + (irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + (irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + 1)))) - ((irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] - 1) - riscv_IRQ_VS_TIMER)] && irq_ctrl_i[(irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + (irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + (irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + 1))) - ((irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] - 1) - riscv_IRQ_VS_TIMER)])
					// Trace: core/decoder.sv:1597:11
					interrupt_cause = INTERRUPTS[interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] - 1)))))-:((interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] - 1)))))) >= (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + 0))))) ? ((interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] - 1)))))) - (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + 0)))))) + 1 : ((interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + 0))))) - (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] - 1))))))) + 1)];
				if (irq_ctrl_i[(irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + (irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + (irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + (irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + 1)))) - ((irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] - 1) - riscv_IRQ_VS_SOFT)] && irq_ctrl_i[(irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + (irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + (irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + 1))) - ((irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] - 1) - riscv_IRQ_VS_SOFT)])
					// Trace: core/decoder.sv:1601:11
					interrupt_cause = INTERRUPTS[interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] - 1))))))))-:((interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] - 1))))))))) >= (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + 0)))))))) ? ((interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] - 1))))))))) - (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + 0))))))))) + 1 : ((interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + 0)))))))) - (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] - 1)))))))))) + 1)];
				if (irq_ctrl_i[(irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + (irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + (irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + (irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + 1)))) - ((irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] - 1) - riscv_IRQ_VS_EXT)] && irq_ctrl_i[(irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + (irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + (irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + 1))) - ((irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] - 1) - riscv_IRQ_VS_EXT)])
					// Trace: core/decoder.sv:1605:11
					interrupt_cause = INTERRUPTS[interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] - 1))-:((interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] - 1))) >= (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + 0)) ? ((interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] - 1))) - (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + 0))) + 1 : ((interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + 0)) - (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] - 1)))) + 1)];
				if (irq_ctrl_i[(irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + (irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + (irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + (irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + 1)))) - ((irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] - 1) - riscv_IRQ_HS_EXT)] && irq_ctrl_i[(irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + (irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + (irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + 1))) - ((irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] - 1) - riscv_IRQ_HS_EXT)])
					// Trace: core/decoder.sv:1609:11
					interrupt_cause = INTERRUPTS[interrupts_t_interrupts_t_CVA6Cfg[17102-:32] - 1-:interrupts_t_interrupts_t_CVA6Cfg[17102-:32]];
			end
			if (CVA6Cfg[16366]) begin
				// Trace: core/decoder.sv:1614:9
				if (irq_ctrl_i[(irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + (irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + (irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + (irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + 1)))) - ((irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] - 1) - riscv_IRQ_S_TIMER)] && irq_ctrl_i[(irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + (irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + (irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + 1))) - ((irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] - 1) - riscv_IRQ_S_TIMER)])
					// Trace: core/decoder.sv:1615:11
					interrupt_cause = INTERRUPTS[interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] - 1))))))-:((interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] - 1))))))) >= (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + 0)))))) ? ((interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] - 1))))))) - (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + 0))))))) + 1 : ((interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + 0)))))) - (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] - 1)))))))) + 1)];
				if (irq_ctrl_i[(irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + (irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + (irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + (irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + 1)))) - ((irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] - 1) - riscv_IRQ_S_SOFT)] && irq_ctrl_i[(irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + (irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + (irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + 1))) - ((irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] - 1) - riscv_IRQ_S_SOFT)])
					// Trace: core/decoder.sv:1619:11
					interrupt_cause = INTERRUPTS[interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] - 1)))))))))-:((interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] - 1)))))))))) >= (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + 0))))))))) ? ((interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] - 1)))))))))) - (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + 0)))))))))) + 1 : ((interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + 0))))))))) - (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] - 1))))))))))) + 1)];
				if (irq_ctrl_i[(irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + (irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + (irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + (irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + 1)))) - ((irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] - 1) - riscv_IRQ_S_EXT)] && (irq_ctrl_i[(irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + (irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + (irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + 1))) - ((irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] - 1) - riscv_IRQ_S_EXT)] | irq_i[ariane_pkg_SupervisorIrq]))
					// Trace: core/decoder.sv:1625:11
					interrupt_cause = INTERRUPTS[interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] - 1)))-:((interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] - 1)))) >= (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + 0))) ? ((interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] - 1)))) - (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + 0)))) + 1 : ((interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + 0))) - (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] - 1))))) + 1)];
			end
			if (irq_ctrl_i[(irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + (irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + (irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + 1))) - ((irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] - 1) - riscv_IRQ_M_TIMER)] && irq_ctrl_i[(irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + (irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + (irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + (irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + 1)))) - ((irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] - 1) - riscv_IRQ_M_TIMER)])
				// Trace: core/decoder.sv:1630:9
				interrupt_cause = INTERRUPTS[interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] - 1))))-:((interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] - 1))))) >= (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + 0)))) ? ((interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] - 1))))) - (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + 0))))) + 1 : ((interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + 0)))) - (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] - 1)))))) + 1)];
			if (irq_ctrl_i[(irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + (irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + (irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + 1))) - ((irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] - 1) - riscv_IRQ_M_SOFT)] && irq_ctrl_i[(irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + (irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + (irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + (irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + 1)))) - ((irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] - 1) - riscv_IRQ_M_SOFT)])
				// Trace: core/decoder.sv:1634:9
				interrupt_cause = INTERRUPTS[interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] - 1)))))))-:((interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] - 1)))))))) >= (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + 0))))))) ? ((interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] - 1)))))))) - (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + 0)))))))) + 1 : ((interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + 0))))))) - (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] - 1))))))))) + 1)];
			if (irq_ctrl_i[(irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + (irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + (irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + 1))) - ((irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] - 1) - riscv_IRQ_M_EXT)] && irq_ctrl_i[(irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + (irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + (irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + (irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + 1)))) - ((irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] - 1) - riscv_IRQ_M_EXT)])
				// Trace: core/decoder.sv:1638:9
				interrupt_cause = INTERRUPTS[interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] - 1)-:((interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] - 1)) >= (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + 0) ? ((interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] - 1)) - (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + 0)) + 1 : ((interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + 0) - (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] + (interrupts_t_interrupts_t_CVA6Cfg[17102-:32] - 1))) + 1)];
			if (interrupt_cause[CVA6Cfg[17102-:32] - 1] && irq_ctrl_i[0]) begin
				begin
					// Trace: core/decoder.sv:1645:9
					if (irq_ctrl_i[(irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + (irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + 1)) - ((irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] - 1) - interrupt_cause[$clog2(CVA6Cfg[17102-:32]) - 1:0])]) begin
						begin
							// Trace: core/decoder.sv:1646:11
							if (CVA6Cfg[16543]) begin : hyp_int_gen
								// Trace: core/decoder.sv:1647:13
								if (v_i && irq_ctrl_i[(irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + 1) - ((irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] - 1) - interrupt_cause[$clog2(CVA6Cfg[17102-:32]) - 1:0])]) begin
									begin
										// Trace: core/decoder.sv:1648:15
										if ((irq_ctrl_i[1] && (priv_lvl_i == 2'b01)) || (priv_lvl_i == 2'b00)) begin
											// Trace: core/decoder.sv:1649:17
											instruction_o[((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) : (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)] = 1'b1;
											// Trace: core/decoder.sv:1650:17
											instruction_o[((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) - ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) : ((((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) + ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) + 1)) - 1)-:((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) + 1)] = interrupt_cause;
										end
									end
								end
								else if (v_i && ~irq_ctrl_i[(irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + 1) - ((irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] - 1) - interrupt_cause[$clog2(CVA6Cfg[17102-:32]) - 1:0])]) begin
									// Trace: core/decoder.sv:1655:15
									instruction_o[((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) : (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)] = 1'b1;
									// Trace: core/decoder.sv:1656:15
									instruction_o[((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) - ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) : ((((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) + ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) + 1)) - 1)-:((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) + 1)] = interrupt_cause;
								end
								else if ((!v_i && ((irq_ctrl_i[1] && (priv_lvl_i == 2'b01)) || (priv_lvl_i == 2'b00))) && ~irq_ctrl_i[(irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] + 1) - ((irq_ctrl_t_irq_ctrl_t_CVA6Cfg[17102-:32] - 1) - interrupt_cause[$clog2(CVA6Cfg[17102-:32]) - 1:0])]) begin
									// Trace: core/decoder.sv:1660:15
									instruction_o[((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) : (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)] = 1'b1;
									// Trace: core/decoder.sv:1661:15
									instruction_o[((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) - ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) : ((((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) + ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) + 1)) - 1)-:((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) + 1)] = interrupt_cause;
								end
							end
							else
								// Trace: core/decoder.sv:1664:13
								if (((CVA6Cfg[16366] && irq_ctrl_i[1]) && (priv_lvl_i == 2'b01)) || (CVA6Cfg[16365] && (priv_lvl_i == 2'b00))) begin
									// Trace: core/decoder.sv:1665:15
									instruction_o[((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) : (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)] = 1'b1;
									// Trace: core/decoder.sv:1666:15
									instruction_o[((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) - ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) : ((((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) + ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) + 1)) - 1)-:((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) + 1)] = interrupt_cause;
								end
						end
					end
					else begin
						// Trace: core/decoder.sv:1670:11
						instruction_o[((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) : (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)] = 1'b1;
						// Trace: core/decoder.sv:1671:11
						instruction_o[((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) - ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) : ((((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) + ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) + 1)) - 1)-:((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) + 1)] = interrupt_cause;
					end
				end
			end
		end
		if ((CVA6Cfg[1321] && debug_req_i) && !debug_mode_i) begin
			// Trace: core/decoder.sv:1678:7
			instruction_o[((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) : (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)] = 1'b1;
			// Trace: core/decoder.sv:1679:7
			instruction_o[((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) - ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) : ((((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) + ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) + 1)) - 1)-:((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) + 1)] = riscv_DEBUG_REQUEST;
		end
	end
	initial _sv2v_0 = 0;
endmodule
