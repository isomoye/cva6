module fpnew_fma_9038D_CD718 (
	clk_i,
	rst_ni,
	operands_i,
	is_boxed_i,
	rnd_mode_i,
	op_i,
	op_mod_i,
	tag_i,
	mask_i,
	aux_i,
	in_valid_i,
	in_ready_o,
	flush_i,
	result_o,
	status_o,
	extension_bit_o,
	tag_o,
	mask_o,
	aux_o,
	out_valid_o,
	out_ready_i,
	busy_o
);
	// removed localparam type TagType_TagType_TagType_TagType_CVA6Cfg_type
	// removed localparam type TagType_TagType_TagType_TagType_config_pkg_NrMaxRules_type
	parameter [17102:0] TagType_TagType_TagType_TagType_CVA6Cfg = 0;
	parameter signed [31:0] TagType_TagType_TagType_TagType_config_pkg_NrMaxRules = 0;
	reg _sv2v_0;
	// Trace: core/cvfpu/src/fpnew_fma.sv:19:13
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	// removed localparam type fpnew_pkg_fp_format_e
	function automatic [2:0] sv2v_cast_5D882;
		input reg [2:0] inp;
		sv2v_cast_5D882 = inp;
	endfunction
	parameter [2:0] FpFormat = sv2v_cast_5D882(0);
	// Trace: core/cvfpu/src/fpnew_fma.sv:20:13
	parameter [31:0] NumPipeRegs = 0;
	// Trace: core/cvfpu/src/fpnew_fma.sv:21:13
	// removed localparam type fpnew_pkg_pipe_config_t
	parameter [1:0] PipeConfig = 2'd0;
	// Trace: core/cvfpu/src/fpnew_fma.sv:22:38
	// removed localparam type TagType
	// Trace: core/cvfpu/src/fpnew_fma.sv:23:38
	// removed localparam type AuxType
	// Trace: core/cvfpu/src/fpnew_fma.sv:25:14
	// removed localparam type fpnew_pkg_fp_encoding_t
	localparam [319:0] fpnew_pkg_FP_ENCODINGS = 320'h8000000170000000b00000034000000050000000a00000005000000020000000800000007;
	function automatic [31:0] fpnew_pkg_fp_width;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:304:44
		input reg [2:0] fmt;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:305:5
		fpnew_pkg_fp_width = (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] + fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32]) + 1;
	endfunction
	localparam [31:0] WIDTH = fpnew_pkg_fp_width(FpFormat);
	// Trace: core/cvfpu/src/fpnew_fma.sv:27:3
	input wire clk_i;
	// Trace: core/cvfpu/src/fpnew_fma.sv:28:3
	input wire rst_ni;
	// Trace: core/cvfpu/src/fpnew_fma.sv:30:3
	input wire [(3 * WIDTH) - 1:0] operands_i;
	// Trace: core/cvfpu/src/fpnew_fma.sv:31:3
	input wire [2:0] is_boxed_i;
	// Trace: core/cvfpu/src/fpnew_fma.sv:32:3
	// removed localparam type fpnew_pkg_roundmode_e
	input wire [2:0] rnd_mode_i;
	// Trace: core/cvfpu/src/fpnew_fma.sv:33:3
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	// removed localparam type fpnew_pkg_operation_e
	input wire [3:0] op_i;
	// Trace: core/cvfpu/src/fpnew_fma.sv:34:3
	input wire op_mod_i;
	// Trace: core/cvfpu/src/fpnew_fma.sv:35:3
	input wire [TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1:0] tag_i;
	// Trace: core/cvfpu/src/fpnew_fma.sv:36:3
	input wire mask_i;
	// Trace: core/cvfpu/src/fpnew_fma.sv:37:3
	input wire aux_i;
	// Trace: core/cvfpu/src/fpnew_fma.sv:39:3
	input wire in_valid_i;
	// Trace: core/cvfpu/src/fpnew_fma.sv:40:3
	output wire in_ready_o;
	// Trace: core/cvfpu/src/fpnew_fma.sv:41:3
	input wire flush_i;
	// Trace: core/cvfpu/src/fpnew_fma.sv:43:3
	output wire [WIDTH - 1:0] result_o;
	// Trace: core/cvfpu/src/fpnew_fma.sv:44:3
	// removed localparam type fpnew_pkg_status_t
	output wire [4:0] status_o;
	// Trace: core/cvfpu/src/fpnew_fma.sv:45:3
	output wire extension_bit_o;
	// Trace: core/cvfpu/src/fpnew_fma.sv:46:3
	output wire [TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1:0] tag_o;
	// Trace: core/cvfpu/src/fpnew_fma.sv:47:3
	output wire mask_o;
	// Trace: core/cvfpu/src/fpnew_fma.sv:48:3
	output wire aux_o;
	// Trace: core/cvfpu/src/fpnew_fma.sv:50:3
	output wire out_valid_o;
	// Trace: core/cvfpu/src/fpnew_fma.sv:51:3
	input wire out_ready_i;
	// Trace: core/cvfpu/src/fpnew_fma.sv:53:3
	output wire busy_o;
	// Trace: core/cvfpu/src/fpnew_fma.sv:59:3
	function automatic [31:0] fpnew_pkg_exp_bits;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:327:44
		input reg [2:0] fmt;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:328:5
		fpnew_pkg_exp_bits = fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32];
	endfunction
	localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(FpFormat);
	// Trace: core/cvfpu/src/fpnew_fma.sv:60:3
	function automatic [31:0] fpnew_pkg_man_bits;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:332:44
		input reg [2:0] fmt;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:333:5
		fpnew_pkg_man_bits = fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32];
	endfunction
	localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(FpFormat);
	// Trace: core/cvfpu/src/fpnew_fma.sv:61:3
	function automatic [31:0] fpnew_pkg_bias;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:337:40
		input reg [2:0] fmt;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:338:5
		fpnew_pkg_bias = $unsigned((2 ** (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] - 1)) - 1);
	endfunction
	localparam [31:0] BIAS = fpnew_pkg_bias(FpFormat);
	// Trace: core/cvfpu/src/fpnew_fma.sv:63:3
	localparam [31:0] PRECISION_BITS = MAN_BITS + 1;
	// Trace: core/cvfpu/src/fpnew_fma.sv:65:3
	localparam [31:0] LOWER_SUM_WIDTH = (2 * PRECISION_BITS) + 3;
	// Trace: core/cvfpu/src/fpnew_fma.sv:66:3
	localparam [31:0] LZC_RESULT_WIDTH = $clog2(LOWER_SUM_WIDTH);
	// Trace: core/cvfpu/src/fpnew_fma.sv:70:3
	function automatic signed [31:0] fpnew_pkg_maximum;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:296:34
		input reg signed [31:0] a;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:296:41
		input reg signed [31:0] b;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:297:5
		fpnew_pkg_maximum = (a > b ? a : b);
	endfunction
	localparam [31:0] EXP_WIDTH = $unsigned(fpnew_pkg_maximum(EXP_BITS + 2, LZC_RESULT_WIDTH));
	// Trace: core/cvfpu/src/fpnew_fma.sv:72:3
	localparam [31:0] SHIFT_AMOUNT_WIDTH = $clog2((3 * PRECISION_BITS) + 5);
	// Trace: core/cvfpu/src/fpnew_fma.sv:74:3
	localparam NUM_INP_REGS = (PipeConfig == 2'd0 ? NumPipeRegs : (PipeConfig == 2'd3 ? (NumPipeRegs + 1) / 3 : 0));
	// Trace: core/cvfpu/src/fpnew_fma.sv:79:3
	localparam NUM_MID_REGS = (PipeConfig == 2'd2 ? NumPipeRegs : (PipeConfig == 2'd3 ? (NumPipeRegs + 2) / 3 : 0));
	// Trace: core/cvfpu/src/fpnew_fma.sv:84:3
	localparam NUM_OUT_REGS = (PipeConfig == 2'd1 ? NumPipeRegs : (PipeConfig == 2'd3 ? NumPipeRegs / 3 : 0));
	// Trace: core/cvfpu/src/fpnew_fma.sv:93:3
	// removed localparam type fp_t
	// Trace: core/cvfpu/src/fpnew_fma.sv:103:3
	reg [((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) - (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0)) + 1) * WIDTH) + (((0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) * WIDTH) - 1) : ((((0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)) + 1) * WIDTH) + (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) * WIDTH) - 1)):((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) * WIDTH : (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) * WIDTH)] inp_pipe_operands_q;
	// Trace: core/cvfpu/src/fpnew_fma.sv:104:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0)] inp_pipe_is_boxed_q;
	// Trace: core/cvfpu/src/fpnew_fma.sv:105:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0)] inp_pipe_rnd_mode_q;
	// Trace: core/cvfpu/src/fpnew_fma.sv:106:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_OP_BITS) + ((NUM_INP_REGS * fpnew_pkg_OP_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_OP_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_OP_BITS : 0)] inp_pipe_op_q;
	// Trace: core/cvfpu/src/fpnew_fma.sv:107:3
	reg [0:NUM_INP_REGS] inp_pipe_op_mod_q;
	// Trace: core/cvfpu/src/fpnew_fma.sv:108:3
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + ((NUM_INP_REGS * TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) - 1) : ((NUM_INP_REGS + 1) * TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] : 0)] inp_pipe_tag_q;
	// Trace: core/cvfpu/src/fpnew_fma.sv:109:3
	reg [0:NUM_INP_REGS] inp_pipe_mask_q;
	// Trace: core/cvfpu/src/fpnew_fma.sv:110:3
	reg [0:NUM_INP_REGS] inp_pipe_aux_q;
	// Trace: core/cvfpu/src/fpnew_fma.sv:111:3
	reg [0:NUM_INP_REGS] inp_pipe_valid_q;
	// Trace: core/cvfpu/src/fpnew_fma.sv:113:3
	wire [0:NUM_INP_REGS] inp_pipe_ready;
	// Trace: core/cvfpu/src/fpnew_fma.sv:116:3
	wire [3 * WIDTH:1] sv2v_tmp_15914;
	assign sv2v_tmp_15914 = operands_i;
	always @(*) inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3 : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3 : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3] = sv2v_tmp_15914;
	// Trace: core/cvfpu/src/fpnew_fma.sv:117:3
	wire [3:1] sv2v_tmp_3D994;
	assign sv2v_tmp_3D994 = is_boxed_i;
	always @(*) inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3+:3] = sv2v_tmp_3D994;
	// Trace: core/cvfpu/src/fpnew_fma.sv:118:3
	wire [3:1] sv2v_tmp_85314;
	assign sv2v_tmp_85314 = rnd_mode_i;
	always @(*) inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3+:3] = sv2v_tmp_85314;
	// Trace: core/cvfpu/src/fpnew_fma.sv:119:3
	wire [4:1] sv2v_tmp_D905E;
	assign sv2v_tmp_D905E = op_i;
	always @(*) inp_pipe_op_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] = sv2v_tmp_D905E;
	// Trace: core/cvfpu/src/fpnew_fma.sv:120:3
	wire [1:1] sv2v_tmp_72E02;
	assign sv2v_tmp_72E02 = op_mod_i;
	always @(*) inp_pipe_op_mod_q[0] = sv2v_tmp_72E02;
	// Trace: core/cvfpu/src/fpnew_fma.sv:121:3
	wire [TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] * 1:1] sv2v_tmp_DE94E;
	assign sv2v_tmp_DE94E = tag_i;
	always @(*) inp_pipe_tag_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]+:TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]] = sv2v_tmp_DE94E;
	// Trace: core/cvfpu/src/fpnew_fma.sv:122:3
	wire [1:1] sv2v_tmp_AE6A6;
	assign sv2v_tmp_AE6A6 = mask_i;
	always @(*) inp_pipe_mask_q[0] = sv2v_tmp_AE6A6;
	// Trace: core/cvfpu/src/fpnew_fma.sv:123:3
	wire [1:1] sv2v_tmp_683C4;
	assign sv2v_tmp_683C4 = aux_i;
	always @(*) inp_pipe_aux_q[0] = sv2v_tmp_683C4;
	// Trace: core/cvfpu/src/fpnew_fma.sv:124:3
	wire [1:1] sv2v_tmp_CFC25;
	assign sv2v_tmp_CFC25 = in_valid_i;
	always @(*) inp_pipe_valid_q[0] = sv2v_tmp_CFC25;
	// Trace: core/cvfpu/src/fpnew_fma.sv:126:3
	assign in_ready_o = inp_pipe_ready[0];
	// Trace: core/cvfpu/src/fpnew_fma.sv:128:3
	genvar _gv_i_66;
	function automatic [3:0] sv2v_cast_4CD2E;
		input reg [3:0] inp;
		sv2v_cast_4CD2E = inp;
	endfunction
	function automatic [TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1:0] sv2v_cast_65D85;
		input reg [TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1:0] inp;
		sv2v_cast_65D85 = inp;
	endfunction
	generate
		for (_gv_i_66 = 0; _gv_i_66 < NUM_INP_REGS; _gv_i_66 = _gv_i_66 + 1) begin : gen_input_pipeline
			localparam i = _gv_i_66;
			// Trace: core/cvfpu/src/fpnew_fma.sv:130:5
			wire reg_ena;
			// Trace: core/cvfpu/src/fpnew_fma.sv:134:5
			assign inp_pipe_ready[i] = inp_pipe_ready[i + 1] | ~inp_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at core/cvfpu/src/fpnew_fma.sv:136:329
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at core/cvfpu/src/fpnew_fma.sv:136:407
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at core/cvfpu/src/fpnew_fma.sv:136:485
					inp_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at core/cvfpu/src/fpnew_fma.sv:136:637
					inp_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (inp_pipe_ready[i] ? inp_pipe_valid_q[i] : inp_pipe_valid_q[i + 1]));
			// Trace: core/cvfpu/src/fpnew_fma.sv:138:5
			assign reg_ena = inp_pipe_ready[i] & inp_pipe_valid_q[i];
			// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:140:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:140:168
				if (!rst_ni)
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:140:265
					inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:140:455
					inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3] <= (reg_ena ? inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3 : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3 : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3] : inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3]);
			// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:141:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:141:168
				if (!rst_ni)
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:141:265
					inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:141:455
					inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= (reg_ena ? inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3+:3] : inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3]);
			// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:142:83
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:142:180
				if (!rst_ni)
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:142:277
					inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:142:467
					inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= (reg_ena ? inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3+:3] : inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3]);
			// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:143:85
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:143:182
				if (!rst_ni)
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:143:279
					inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= sv2v_cast_4CD2E(0);
				else
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:143:469
					inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= (reg_ena ? inp_pipe_op_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] : inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS]);
			// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:144:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:144:168
				if (!rst_ni)
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:144:265
					inp_pipe_op_mod_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:144:455
					inp_pipe_op_mod_q[i + 1] <= (reg_ena ? inp_pipe_op_mod_q[i] : inp_pipe_op_mod_q[i + 1]);
			// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:145:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:145:178
				if (!rst_ni)
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:145:275
					inp_pipe_tag_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]+:TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]] <= sv2v_cast_65D85(1'sb0);
				else
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:145:465
					inp_pipe_tag_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]+:TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]] <= (reg_ena ? inp_pipe_tag_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]+:TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]] : inp_pipe_tag_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]+:TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]]);
			// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:146:71
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:146:168
				if (!rst_ni)
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:146:265
					inp_pipe_mask_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:146:455
					inp_pipe_mask_q[i + 1] <= (reg_ena ? inp_pipe_mask_q[i] : inp_pipe_mask_q[i + 1]);
			// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:147:81
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:147:178
				if (!rst_ni)
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:147:275
					inp_pipe_aux_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:147:465
					inp_pipe_aux_q[i + 1] <= (reg_ena ? inp_pipe_aux_q[i] : inp_pipe_aux_q[i + 1]);
		end
	endgenerate
	// Trace: core/cvfpu/src/fpnew_fma.sv:153:3
	// removed localparam type fpnew_pkg_fp_info_t
	wire [23:0] info_q;
	// Trace: core/cvfpu/src/fpnew_fma.sv:156:3
	fpnew_classifier #(
		.FpFormat(FpFormat),
		.NumOperands(3)
	) i_class_inputs(
		.operands_i(inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3 : ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3 : ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3]),
		.is_boxed_i(inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3]),
		.info_o(info_q)
	);
	// Trace: core/cvfpu/src/fpnew_fma.sv:165:3
	reg [((1 + EXP_BITS) + MAN_BITS) - 1:0] operand_a;
	reg [((1 + EXP_BITS) + MAN_BITS) - 1:0] operand_b;
	reg [((1 + EXP_BITS) + MAN_BITS) - 1:0] operand_c;
	// Trace: core/cvfpu/src/fpnew_fma.sv:166:3
	reg [7:0] info_a;
	reg [7:0] info_b;
	reg [7:0] info_c;
	// Trace: core/cvfpu/src/fpnew_fma.sv:180:3
	localparam [0:0] fpnew_pkg_DONT_CARE = 1'b1;
	function automatic [EXP_BITS - 1:0] sv2v_cast_51E93;
		input reg [EXP_BITS - 1:0] inp;
		sv2v_cast_51E93 = inp;
	endfunction
	function automatic [MAN_BITS - 1:0] sv2v_cast_78D38;
		input reg [MAN_BITS - 1:0] inp;
		sv2v_cast_78D38 = inp;
	endfunction
	function automatic [EXP_BITS - 1:0] sv2v_cast_89227;
		input reg [EXP_BITS - 1:0] inp;
		sv2v_cast_89227 = inp;
	endfunction
	function automatic [MAN_BITS - 1:0] sv2v_cast_D5F4C;
		input reg [MAN_BITS - 1:0] inp;
		sv2v_cast_D5F4C = inp;
	endfunction
	always @(*) begin : op_select
		if (_sv2v_0)
			;
		// Trace: core/cvfpu/src/fpnew_fma.sv:183:5
		operand_a = inp_pipe_operands_q[((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3 : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1))) * WIDTH+:WIDTH];
		// Trace: core/cvfpu/src/fpnew_fma.sv:184:5
		operand_b = inp_pipe_operands_q[((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3) + 1 : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - ((((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1))) * WIDTH+:WIDTH];
		// Trace: core/cvfpu/src/fpnew_fma.sv:185:5
		operand_c = inp_pipe_operands_q[((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3) + 2 : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - ((((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1))) * WIDTH+:WIDTH];
		// Trace: core/cvfpu/src/fpnew_fma.sv:186:5
		info_a = info_q[0+:8];
		// Trace: core/cvfpu/src/fpnew_fma.sv:187:5
		info_b = info_q[8+:8];
		// Trace: core/cvfpu/src/fpnew_fma.sv:188:5
		info_c = info_q[16+:8];
		// Trace: core/cvfpu/src/fpnew_fma.sv:191:5
		operand_c[1 + (EXP_BITS + (MAN_BITS - 1))] = operand_c[1 + (EXP_BITS + (MAN_BITS - 1))] ^ inp_pipe_op_mod_q[NUM_INP_REGS];
		// Trace: core/cvfpu/src/fpnew_fma.sv:193:5
		(* full_case, parallel_case *)
		case (inp_pipe_op_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS])
			sv2v_cast_4CD2E(0):
				;
			sv2v_cast_4CD2E(1):
				// Trace: core/cvfpu/src/fpnew_fma.sv:195:26
				operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] = ~operand_a[1 + (EXP_BITS + (MAN_BITS - 1))];
			sv2v_cast_4CD2E(2): begin
				// Trace: core/cvfpu/src/fpnew_fma.sv:197:9
				operand_a = {1'b0, sv2v_cast_51E93(BIAS), sv2v_cast_78D38(1'sb0)};
				// Trace: core/cvfpu/src/fpnew_fma.sv:198:9
				info_a = 8'b10000001;
			end
			sv2v_cast_4CD2E(3): begin
				// Trace: core/cvfpu/src/fpnew_fma.sv:201:9
				if (inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3] == 3'b010)
					// Trace: core/cvfpu/src/fpnew_fma.sv:202:11
					operand_c = {1'b0, sv2v_cast_89227(1'sb0), sv2v_cast_78D38(1'sb0)};
				else
					// Trace: core/cvfpu/src/fpnew_fma.sv:204:11
					operand_c = {1'b1, sv2v_cast_89227(1'sb0), sv2v_cast_78D38(1'sb0)};
				// Trace: core/cvfpu/src/fpnew_fma.sv:205:9
				info_c = 8'b00100001;
			end
			default: begin
				// Trace: core/cvfpu/src/fpnew_fma.sv:208:9
				operand_a = {fpnew_pkg_DONT_CARE, sv2v_cast_51E93(fpnew_pkg_DONT_CARE), sv2v_cast_D5F4C(fpnew_pkg_DONT_CARE)};
				// Trace: core/cvfpu/src/fpnew_fma.sv:209:9
				operand_b = {fpnew_pkg_DONT_CARE, sv2v_cast_51E93(fpnew_pkg_DONT_CARE), sv2v_cast_D5F4C(fpnew_pkg_DONT_CARE)};
				// Trace: core/cvfpu/src/fpnew_fma.sv:210:9
				operand_c = {fpnew_pkg_DONT_CARE, sv2v_cast_51E93(fpnew_pkg_DONT_CARE), sv2v_cast_D5F4C(fpnew_pkg_DONT_CARE)};
				// Trace: core/cvfpu/src/fpnew_fma.sv:211:9
				info_a = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
				// Trace: core/cvfpu/src/fpnew_fma.sv:212:9
				info_b = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
				// Trace: core/cvfpu/src/fpnew_fma.sv:213:9
				info_c = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
			end
		endcase
	end
	// Trace: core/cvfpu/src/fpnew_fma.sv:221:3
	wire any_operand_inf;
	// Trace: core/cvfpu/src/fpnew_fma.sv:222:3
	wire any_operand_nan;
	// Trace: core/cvfpu/src/fpnew_fma.sv:223:3
	wire signalling_nan;
	// Trace: core/cvfpu/src/fpnew_fma.sv:224:3
	wire effective_subtraction;
	// Trace: core/cvfpu/src/fpnew_fma.sv:225:3
	wire tentative_sign;
	// Trace: core/cvfpu/src/fpnew_fma.sv:228:3
	assign any_operand_inf = |{info_a[4], info_b[4], info_c[4]};
	// Trace: core/cvfpu/src/fpnew_fma.sv:229:3
	assign any_operand_nan = |{info_a[3], info_b[3], info_c[3]};
	// Trace: core/cvfpu/src/fpnew_fma.sv:230:3
	assign signalling_nan = |{info_a[2], info_b[2], info_c[2]};
	// Trace: core/cvfpu/src/fpnew_fma.sv:232:3
	assign effective_subtraction = (operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] ^ operand_b[1 + (EXP_BITS + (MAN_BITS - 1))]) ^ operand_c[1 + (EXP_BITS + (MAN_BITS - 1))];
	// Trace: core/cvfpu/src/fpnew_fma.sv:234:3
	assign tentative_sign = operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] ^ operand_b[1 + (EXP_BITS + (MAN_BITS - 1))];
	// Trace: core/cvfpu/src/fpnew_fma.sv:239:3
	reg [((1 + EXP_BITS) + MAN_BITS) - 1:0] special_result;
	// Trace: core/cvfpu/src/fpnew_fma.sv:240:3
	reg [4:0] special_status;
	// Trace: core/cvfpu/src/fpnew_fma.sv:241:3
	reg result_is_special;
	// Trace: core/cvfpu/src/fpnew_fma.sv:243:3
	always @(*) begin : special_cases
		if (_sv2v_0)
			;
		// Trace: core/cvfpu/src/fpnew_fma.sv:245:5
		special_result = {1'b0, sv2v_cast_89227(1'sb1), sv2v_cast_D5F4C(2 ** (MAN_BITS - 1))};
		// Trace: core/cvfpu/src/fpnew_fma.sv:246:5
		special_status = 1'sb0;
		// Trace: core/cvfpu/src/fpnew_fma.sv:247:5
		result_is_special = 1'b0;
		// Trace: core/cvfpu/src/fpnew_fma.sv:253:5
		if ((info_a[4] && info_b[5]) || (info_a[5] && info_b[4])) begin
			// Trace: core/cvfpu/src/fpnew_fma.sv:254:7
			result_is_special = 1'b1;
			// Trace: core/cvfpu/src/fpnew_fma.sv:255:7
			special_status[4] = 1'b1;
		end
		else if (any_operand_nan) begin
			// Trace: core/cvfpu/src/fpnew_fma.sv:258:7
			result_is_special = 1'b1;
			// Trace: core/cvfpu/src/fpnew_fma.sv:259:7
			special_status[4] = signalling_nan;
		end
		else if (any_operand_inf) begin
			// Trace: core/cvfpu/src/fpnew_fma.sv:262:7
			result_is_special = 1'b1;
			// Trace: core/cvfpu/src/fpnew_fma.sv:264:7
			if (((info_a[4] || info_b[4]) && info_c[4]) && effective_subtraction)
				// Trace: core/cvfpu/src/fpnew_fma.sv:265:9
				special_status[4] = 1'b1;
			else if (info_a[4] || info_b[4])
				// Trace: core/cvfpu/src/fpnew_fma.sv:269:9
				special_result = {operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] ^ operand_b[1 + (EXP_BITS + (MAN_BITS - 1))], sv2v_cast_89227(1'sb1), sv2v_cast_78D38(1'sb0)};
			else if (info_c[4])
				// Trace: core/cvfpu/src/fpnew_fma.sv:273:9
				special_result = {operand_c[1 + (EXP_BITS + (MAN_BITS - 1))], sv2v_cast_89227(1'sb1), sv2v_cast_78D38(1'sb0)};
		end
	end
	// Trace: core/cvfpu/src/fpnew_fma.sv:281:3
	wire signed [EXP_WIDTH - 1:0] exponent_a;
	wire signed [EXP_WIDTH - 1:0] exponent_b;
	wire signed [EXP_WIDTH - 1:0] exponent_c;
	// Trace: core/cvfpu/src/fpnew_fma.sv:282:3
	wire signed [EXP_WIDTH - 1:0] exponent_addend;
	wire signed [EXP_WIDTH - 1:0] exponent_product;
	wire signed [EXP_WIDTH - 1:0] exponent_difference;
	// Trace: core/cvfpu/src/fpnew_fma.sv:283:3
	wire signed [EXP_WIDTH - 1:0] tentative_exponent;
	// Trace: core/cvfpu/src/fpnew_fma.sv:286:3
	assign exponent_a = $signed({1'b0, operand_a[EXP_BITS + (MAN_BITS - 1)-:((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1)]});
	// Trace: core/cvfpu/src/fpnew_fma.sv:287:3
	assign exponent_b = $signed({1'b0, operand_b[EXP_BITS + (MAN_BITS - 1)-:((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1)]});
	// Trace: core/cvfpu/src/fpnew_fma.sv:288:3
	assign exponent_c = $signed({1'b0, operand_c[EXP_BITS + (MAN_BITS - 1)-:((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1)]});
	// Trace: core/cvfpu/src/fpnew_fma.sv:292:3
	assign exponent_addend = $signed(exponent_c + $signed({1'b0, ~info_c[7]}));
	// Trace: core/cvfpu/src/fpnew_fma.sv:294:3
	assign exponent_product = (info_a[5] || info_b[5] ? 2 - $signed(BIAS) : $signed((((exponent_a + info_a[6]) + exponent_b) + info_b[6]) - $signed(BIAS)));
	// Trace: core/cvfpu/src/fpnew_fma.sv:300:3
	assign exponent_difference = exponent_addend - exponent_product;
	// Trace: core/cvfpu/src/fpnew_fma.sv:302:3
	assign tentative_exponent = (exponent_difference > 0 ? exponent_addend : exponent_product);
	// Trace: core/cvfpu/src/fpnew_fma.sv:305:3
	reg [SHIFT_AMOUNT_WIDTH - 1:0] addend_shamt;
	// Trace: core/cvfpu/src/fpnew_fma.sv:307:3
	always @(*) begin : addend_shift_amount
		if (_sv2v_0)
			;
		// Trace: core/cvfpu/src/fpnew_fma.sv:309:5
		if (exponent_difference <= $signed((-2 * PRECISION_BITS) - 1))
			// Trace: core/cvfpu/src/fpnew_fma.sv:310:7
			addend_shamt = (3 * PRECISION_BITS) + 4;
		else if (exponent_difference <= $signed(PRECISION_BITS + 2))
			// Trace: core/cvfpu/src/fpnew_fma.sv:313:7
			addend_shamt = $unsigned(($signed(PRECISION_BITS) + 3) - exponent_difference);
		else
			// Trace: core/cvfpu/src/fpnew_fma.sv:316:7
			addend_shamt = 0;
	end
	// Trace: core/cvfpu/src/fpnew_fma.sv:322:3
	wire [PRECISION_BITS - 1:0] mantissa_a;
	wire [PRECISION_BITS - 1:0] mantissa_b;
	wire [PRECISION_BITS - 1:0] mantissa_c;
	// Trace: core/cvfpu/src/fpnew_fma.sv:323:3
	wire [(2 * PRECISION_BITS) - 1:0] product;
	// Trace: core/cvfpu/src/fpnew_fma.sv:324:3
	wire [(3 * PRECISION_BITS) + 3:0] product_shifted;
	// Trace: core/cvfpu/src/fpnew_fma.sv:327:3
	assign mantissa_a = {info_a[7], operand_a[MAN_BITS - 1-:MAN_BITS]};
	// Trace: core/cvfpu/src/fpnew_fma.sv:328:3
	assign mantissa_b = {info_b[7], operand_b[MAN_BITS - 1-:MAN_BITS]};
	// Trace: core/cvfpu/src/fpnew_fma.sv:329:3
	assign mantissa_c = {info_c[7], operand_c[MAN_BITS - 1-:MAN_BITS]};
	// Trace: core/cvfpu/src/fpnew_fma.sv:332:3
	assign product = mantissa_a * mantissa_b;
	// Trace: core/cvfpu/src/fpnew_fma.sv:337:3
	assign product_shifted = product << 2;
	// Trace: core/cvfpu/src/fpnew_fma.sv:342:3
	wire [(3 * PRECISION_BITS) + 3:0] addend_after_shift;
	// Trace: core/cvfpu/src/fpnew_fma.sv:343:3
	wire [PRECISION_BITS - 1:0] addend_sticky_bits;
	// Trace: core/cvfpu/src/fpnew_fma.sv:344:3
	wire sticky_before_add;
	// Trace: core/cvfpu/src/fpnew_fma.sv:345:3
	wire [(3 * PRECISION_BITS) + 3:0] addend_shifted;
	// Trace: core/cvfpu/src/fpnew_fma.sv:346:3
	wire inject_carry_in;
	// Trace: core/cvfpu/src/fpnew_fma.sv:356:3
	assign {addend_after_shift, addend_sticky_bits} = (mantissa_c << ((3 * PRECISION_BITS) + 4)) >> addend_shamt;
	// Trace: core/cvfpu/src/fpnew_fma.sv:359:3
	assign sticky_before_add = |addend_sticky_bits;
	// Trace: core/cvfpu/src/fpnew_fma.sv:363:3
	assign addend_shifted = (effective_subtraction ? ~addend_after_shift : addend_after_shift);
	// Trace: core/cvfpu/src/fpnew_fma.sv:364:3
	assign inject_carry_in = effective_subtraction & ~sticky_before_add;
	// Trace: core/cvfpu/src/fpnew_fma.sv:369:3
	wire [(3 * PRECISION_BITS) + 4:0] sum_raw;
	// Trace: core/cvfpu/src/fpnew_fma.sv:370:3
	wire sum_carry;
	// Trace: core/cvfpu/src/fpnew_fma.sv:371:3
	wire [(3 * PRECISION_BITS) + 3:0] sum;
	// Trace: core/cvfpu/src/fpnew_fma.sv:372:3
	wire final_sign;
	// Trace: core/cvfpu/src/fpnew_fma.sv:375:3
	assign sum_raw = (product_shifted + addend_shifted) + inject_carry_in;
	// Trace: core/cvfpu/src/fpnew_fma.sv:376:3
	assign sum_carry = sum_raw[(3 * PRECISION_BITS) + 4];
	// Trace: core/cvfpu/src/fpnew_fma.sv:379:3
	assign sum = (effective_subtraction && ~sum_carry ? -sum_raw : sum_raw);
	// Trace: core/cvfpu/src/fpnew_fma.sv:382:3
	assign final_sign = (effective_subtraction && (sum_carry == tentative_sign) ? 1'b1 : (effective_subtraction ? 1'b0 : tentative_sign));
	// Trace: core/cvfpu/src/fpnew_fma.sv:390:3
	wire effective_subtraction_q;
	// Trace: core/cvfpu/src/fpnew_fma.sv:391:3
	wire signed [EXP_WIDTH - 1:0] exponent_product_q;
	// Trace: core/cvfpu/src/fpnew_fma.sv:392:3
	wire signed [EXP_WIDTH - 1:0] exponent_difference_q;
	// Trace: core/cvfpu/src/fpnew_fma.sv:393:3
	wire signed [EXP_WIDTH - 1:0] tentative_exponent_q;
	// Trace: core/cvfpu/src/fpnew_fma.sv:394:3
	wire [SHIFT_AMOUNT_WIDTH - 1:0] addend_shamt_q;
	// Trace: core/cvfpu/src/fpnew_fma.sv:395:3
	wire sticky_before_add_q;
	// Trace: core/cvfpu/src/fpnew_fma.sv:396:3
	wire [(3 * PRECISION_BITS) + 3:0] sum_q;
	// Trace: core/cvfpu/src/fpnew_fma.sv:397:3
	wire final_sign_q;
	// Trace: core/cvfpu/src/fpnew_fma.sv:398:3
	wire [2:0] rnd_mode_q;
	// Trace: core/cvfpu/src/fpnew_fma.sv:399:3
	wire result_is_special_q;
	// Trace: core/cvfpu/src/fpnew_fma.sv:400:3
	wire [((1 + EXP_BITS) + MAN_BITS) - 1:0] special_result_q;
	// Trace: core/cvfpu/src/fpnew_fma.sv:401:3
	wire [4:0] special_status_q;
	// Trace: core/cvfpu/src/fpnew_fma.sv:403:3
	reg [0:NUM_MID_REGS] mid_pipe_eff_sub_q;
	// Trace: core/cvfpu/src/fpnew_fma.sv:404:3
	reg signed [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * EXP_WIDTH) + ((NUM_MID_REGS * EXP_WIDTH) - 1) : ((NUM_MID_REGS + 1) * EXP_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * EXP_WIDTH : 0)] mid_pipe_exp_prod_q;
	// Trace: core/cvfpu/src/fpnew_fma.sv:405:3
	reg signed [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * EXP_WIDTH) + ((NUM_MID_REGS * EXP_WIDTH) - 1) : ((NUM_MID_REGS + 1) * EXP_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * EXP_WIDTH : 0)] mid_pipe_exp_diff_q;
	// Trace: core/cvfpu/src/fpnew_fma.sv:406:3
	reg signed [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * EXP_WIDTH) + ((NUM_MID_REGS * EXP_WIDTH) - 1) : ((NUM_MID_REGS + 1) * EXP_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * EXP_WIDTH : 0)] mid_pipe_tent_exp_q;
	// Trace: core/cvfpu/src/fpnew_fma.sv:407:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * SHIFT_AMOUNT_WIDTH) + ((NUM_MID_REGS * SHIFT_AMOUNT_WIDTH) - 1) : ((NUM_MID_REGS + 1) * SHIFT_AMOUNT_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * SHIFT_AMOUNT_WIDTH : 0)] mid_pipe_add_shamt_q;
	// Trace: core/cvfpu/src/fpnew_fma.sv:408:3
	reg [0:NUM_MID_REGS] mid_pipe_sticky_q;
	// Trace: core/cvfpu/src/fpnew_fma.sv:409:3
	reg [(0 >= NUM_MID_REGS ? (((3 * PRECISION_BITS) + 3) >= 0 ? ((1 - NUM_MID_REGS) * ((3 * PRECISION_BITS) + 4)) + ((NUM_MID_REGS * ((3 * PRECISION_BITS) + 4)) - 1) : ((1 - NUM_MID_REGS) * (1 - ((3 * PRECISION_BITS) + 3))) + ((((3 * PRECISION_BITS) + 3) + (NUM_MID_REGS * (1 - ((3 * PRECISION_BITS) + 3)))) - 1)) : (((3 * PRECISION_BITS) + 3) >= 0 ? ((NUM_MID_REGS + 1) * ((3 * PRECISION_BITS) + 4)) - 1 : ((NUM_MID_REGS + 1) * (1 - ((3 * PRECISION_BITS) + 3))) + ((3 * PRECISION_BITS) + 2))):(0 >= NUM_MID_REGS ? (((3 * PRECISION_BITS) + 3) >= 0 ? NUM_MID_REGS * ((3 * PRECISION_BITS) + 4) : ((3 * PRECISION_BITS) + 3) + (NUM_MID_REGS * (1 - ((3 * PRECISION_BITS) + 3)))) : (((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3))] mid_pipe_sum_q;
	// Trace: core/cvfpu/src/fpnew_fma.sv:410:3
	reg [0:NUM_MID_REGS] mid_pipe_final_sign_q;
	// Trace: core/cvfpu/src/fpnew_fma.sv:411:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * 3) + ((NUM_MID_REGS * 3) - 1) : ((NUM_MID_REGS + 1) * 3) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * 3 : 0)] mid_pipe_rnd_mode_q;
	// Trace: core/cvfpu/src/fpnew_fma.sv:412:3
	reg [0:NUM_MID_REGS] mid_pipe_res_is_spec_q;
	// Trace: core/cvfpu/src/fpnew_fma.sv:413:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * ((1 + EXP_BITS) + MAN_BITS)) + ((NUM_MID_REGS * ((1 + EXP_BITS) + MAN_BITS)) - 1) : ((NUM_MID_REGS + 1) * ((1 + EXP_BITS) + MAN_BITS)) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * ((1 + EXP_BITS) + MAN_BITS) : 0)] mid_pipe_spec_res_q;
	// Trace: core/cvfpu/src/fpnew_fma.sv:414:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * 5) + ((NUM_MID_REGS * 5) - 1) : ((NUM_MID_REGS + 1) * 5) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * 5 : 0)] mid_pipe_spec_stat_q;
	// Trace: core/cvfpu/src/fpnew_fma.sv:415:3
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + ((NUM_MID_REGS * TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) - 1) : ((NUM_MID_REGS + 1) * TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] : 0)] mid_pipe_tag_q;
	// Trace: core/cvfpu/src/fpnew_fma.sv:416:3
	reg [0:NUM_MID_REGS] mid_pipe_mask_q;
	// Trace: core/cvfpu/src/fpnew_fma.sv:417:3
	reg [0:NUM_MID_REGS] mid_pipe_aux_q;
	// Trace: core/cvfpu/src/fpnew_fma.sv:418:3
	reg [0:NUM_MID_REGS] mid_pipe_valid_q;
	// Trace: core/cvfpu/src/fpnew_fma.sv:420:3
	wire [0:NUM_MID_REGS] mid_pipe_ready;
	// Trace: core/cvfpu/src/fpnew_fma.sv:423:3
	wire [1:1] sv2v_tmp_301F1;
	assign sv2v_tmp_301F1 = effective_subtraction;
	always @(*) mid_pipe_eff_sub_q[0] = sv2v_tmp_301F1;
	// Trace: core/cvfpu/src/fpnew_fma.sv:424:3
	wire [EXP_WIDTH * 1:1] sv2v_tmp_27C8D;
	assign sv2v_tmp_27C8D = exponent_product;
	always @(*) mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH] = sv2v_tmp_27C8D;
	// Trace: core/cvfpu/src/fpnew_fma.sv:425:3
	wire [EXP_WIDTH * 1:1] sv2v_tmp_DEAE0;
	assign sv2v_tmp_DEAE0 = exponent_difference;
	always @(*) mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH] = sv2v_tmp_DEAE0;
	// Trace: core/cvfpu/src/fpnew_fma.sv:426:3
	wire [EXP_WIDTH * 1:1] sv2v_tmp_530A2;
	assign sv2v_tmp_530A2 = tentative_exponent;
	always @(*) mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH] = sv2v_tmp_530A2;
	// Trace: core/cvfpu/src/fpnew_fma.sv:427:3
	wire [SHIFT_AMOUNT_WIDTH * 1:1] sv2v_tmp_12F7F;
	assign sv2v_tmp_12F7F = addend_shamt;
	always @(*) mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH] = sv2v_tmp_12F7F;
	// Trace: core/cvfpu/src/fpnew_fma.sv:428:3
	wire [1:1] sv2v_tmp_6A24C;
	assign sv2v_tmp_6A24C = sticky_before_add;
	always @(*) mid_pipe_sticky_q[0] = sv2v_tmp_6A24C;
	// Trace: core/cvfpu/src/fpnew_fma.sv:429:3
	wire [(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)) * 1:1] sv2v_tmp_A48E2;
	assign sv2v_tmp_A48E2 = sum;
	always @(*) mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))] = sv2v_tmp_A48E2;
	// Trace: core/cvfpu/src/fpnew_fma.sv:430:3
	wire [1:1] sv2v_tmp_9C379;
	assign sv2v_tmp_9C379 = final_sign;
	always @(*) mid_pipe_final_sign_q[0] = sv2v_tmp_9C379;
	// Trace: core/cvfpu/src/fpnew_fma.sv:431:3
	wire [3:1] sv2v_tmp_C990F;
	assign sv2v_tmp_C990F = inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3];
	always @(*) mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * 3+:3] = sv2v_tmp_C990F;
	// Trace: core/cvfpu/src/fpnew_fma.sv:432:3
	wire [1:1] sv2v_tmp_08378;
	assign sv2v_tmp_08378 = result_is_special;
	always @(*) mid_pipe_res_is_spec_q[0] = sv2v_tmp_08378;
	// Trace: core/cvfpu/src/fpnew_fma.sv:433:3
	wire [((1 + EXP_BITS) + MAN_BITS) * 1:1] sv2v_tmp_8913F;
	assign sv2v_tmp_8913F = special_result;
	always @(*) mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] = sv2v_tmp_8913F;
	// Trace: core/cvfpu/src/fpnew_fma.sv:434:3
	wire [5:1] sv2v_tmp_9D338;
	assign sv2v_tmp_9D338 = special_status;
	always @(*) mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * 5+:5] = sv2v_tmp_9D338;
	// Trace: core/cvfpu/src/fpnew_fma.sv:435:3
	wire [TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] * 1:1] sv2v_tmp_339B9;
	assign sv2v_tmp_339B9 = inp_pipe_tag_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]+:TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]];
	always @(*) mid_pipe_tag_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]+:TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]] = sv2v_tmp_339B9;
	// Trace: core/cvfpu/src/fpnew_fma.sv:436:3
	wire [1:1] sv2v_tmp_FAFEF;
	assign sv2v_tmp_FAFEF = inp_pipe_mask_q[NUM_INP_REGS];
	always @(*) mid_pipe_mask_q[0] = sv2v_tmp_FAFEF;
	// Trace: core/cvfpu/src/fpnew_fma.sv:437:3
	wire [1:1] sv2v_tmp_8CE3D;
	assign sv2v_tmp_8CE3D = inp_pipe_aux_q[NUM_INP_REGS];
	always @(*) mid_pipe_aux_q[0] = sv2v_tmp_8CE3D;
	// Trace: core/cvfpu/src/fpnew_fma.sv:438:3
	wire [1:1] sv2v_tmp_C7159;
	assign sv2v_tmp_C7159 = inp_pipe_valid_q[NUM_INP_REGS];
	always @(*) mid_pipe_valid_q[0] = sv2v_tmp_C7159;
	// Trace: core/cvfpu/src/fpnew_fma.sv:440:3
	assign inp_pipe_ready[NUM_INP_REGS] = mid_pipe_ready[0];
	// Trace: core/cvfpu/src/fpnew_fma.sv:443:3
	genvar _gv_i_67;
	generate
		for (_gv_i_67 = 0; _gv_i_67 < NUM_MID_REGS; _gv_i_67 = _gv_i_67 + 1) begin : gen_inside_pipeline
			localparam i = _gv_i_67;
			// Trace: core/cvfpu/src/fpnew_fma.sv:445:5
			wire reg_ena;
			// Trace: core/cvfpu/src/fpnew_fma.sv:449:5
			assign mid_pipe_ready[i] = mid_pipe_ready[i + 1] | ~mid_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at core/cvfpu/src/fpnew_fma.sv:451:329
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at core/cvfpu/src/fpnew_fma.sv:451:407
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at core/cvfpu/src/fpnew_fma.sv:451:485
					mid_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at core/cvfpu/src/fpnew_fma.sv:451:637
					mid_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (mid_pipe_ready[i] ? mid_pipe_valid_q[i] : mid_pipe_valid_q[i + 1]));
			// Trace: core/cvfpu/src/fpnew_fma.sv:453:5
			assign reg_ena = mid_pipe_ready[i] & mid_pipe_valid_q[i];
			// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:455:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:455:174
				if (!rst_ni)
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:455:271
					mid_pipe_eff_sub_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:455:461
					mid_pipe_eff_sub_q[i + 1] <= (reg_ena ? mid_pipe_eff_sub_q[i] : mid_pipe_eff_sub_q[i + 1]);
			// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:456:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:456:174
				if (!rst_ni)
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:456:271
					mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:456:461
					mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= (reg_ena ? mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * EXP_WIDTH+:EXP_WIDTH] : mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH]);
			// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:457:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:457:174
				if (!rst_ni)
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:457:271
					mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:457:461
					mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= (reg_ena ? mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * EXP_WIDTH+:EXP_WIDTH] : mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH]);
			// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:458:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:458:174
				if (!rst_ni)
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:458:271
					mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:458:461
					mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= (reg_ena ? mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * EXP_WIDTH+:EXP_WIDTH] : mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH]);
			// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:459:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:459:174
				if (!rst_ni)
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:459:271
					mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:459:461
					mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH] <= (reg_ena ? mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH] : mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH]);
			// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:460:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:460:174
				if (!rst_ni)
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:460:271
					mid_pipe_sticky_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:460:461
					mid_pipe_sticky_q[i + 1] <= (reg_ena ? mid_pipe_sticky_q[i] : mid_pipe_sticky_q[i + 1]);
			// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:461:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:461:174
				if (!rst_ni)
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:461:271
					mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:461:461
					mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))] <= (reg_ena ? mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))] : mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))]);
			// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:462:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:462:174
				if (!rst_ni)
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:462:271
					mid_pipe_final_sign_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:462:461
					mid_pipe_final_sign_q[i + 1] <= (reg_ena ? mid_pipe_final_sign_q[i] : mid_pipe_final_sign_q[i + 1]);
			// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:463:89
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:463:186
				if (!rst_ni)
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:463:283
					mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:463:473
					mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3] <= (reg_ena ? mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * 3+:3] : mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3]);
			// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:464:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:464:174
				if (!rst_ni)
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:464:271
					mid_pipe_res_is_spec_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:464:461
					mid_pipe_res_is_spec_q[i + 1] <= (reg_ena ? mid_pipe_res_is_spec_q[i] : mid_pipe_res_is_spec_q[i + 1]);
			// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:465:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:465:174
				if (!rst_ni)
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:465:271
					mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:465:461
					mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] <= (reg_ena ? mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] : mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS]);
			// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:466:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:466:174
				if (!rst_ni)
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:466:271
					mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 5+:5] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:466:461
					mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 5+:5] <= (reg_ena ? mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * 5+:5] : mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 5+:5]);
			// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:467:87
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:467:184
				if (!rst_ni)
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:467:281
					mid_pipe_tag_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]+:TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]] <= sv2v_cast_65D85(1'sb0);
				else
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:467:471
					mid_pipe_tag_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]+:TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]] <= (reg_ena ? mid_pipe_tag_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]+:TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]] : mid_pipe_tag_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]+:TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]]);
			// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:468:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:468:174
				if (!rst_ni)
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:468:271
					mid_pipe_mask_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:468:461
					mid_pipe_mask_q[i + 1] <= (reg_ena ? mid_pipe_mask_q[i] : mid_pipe_mask_q[i + 1]);
			// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:469:87
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:469:184
				if (!rst_ni)
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:469:281
					mid_pipe_aux_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:469:471
					mid_pipe_aux_q[i + 1] <= (reg_ena ? mid_pipe_aux_q[i] : mid_pipe_aux_q[i + 1]);
		end
	endgenerate
	// Trace: core/cvfpu/src/fpnew_fma.sv:472:3
	assign effective_subtraction_q = mid_pipe_eff_sub_q[NUM_MID_REGS];
	// Trace: core/cvfpu/src/fpnew_fma.sv:473:3
	assign exponent_product_q = mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH];
	// Trace: core/cvfpu/src/fpnew_fma.sv:474:3
	assign exponent_difference_q = mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH];
	// Trace: core/cvfpu/src/fpnew_fma.sv:475:3
	assign tentative_exponent_q = mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH];
	// Trace: core/cvfpu/src/fpnew_fma.sv:476:3
	assign addend_shamt_q = mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH];
	// Trace: core/cvfpu/src/fpnew_fma.sv:477:3
	assign sticky_before_add_q = mid_pipe_sticky_q[NUM_MID_REGS];
	// Trace: core/cvfpu/src/fpnew_fma.sv:478:3
	assign sum_q = mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))];
	// Trace: core/cvfpu/src/fpnew_fma.sv:479:3
	assign final_sign_q = mid_pipe_final_sign_q[NUM_MID_REGS];
	// Trace: core/cvfpu/src/fpnew_fma.sv:480:3
	assign rnd_mode_q = mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * 3+:3];
	// Trace: core/cvfpu/src/fpnew_fma.sv:481:3
	assign result_is_special_q = mid_pipe_res_is_spec_q[NUM_MID_REGS];
	// Trace: core/cvfpu/src/fpnew_fma.sv:482:3
	assign special_result_q = mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS];
	// Trace: core/cvfpu/src/fpnew_fma.sv:483:3
	assign special_status_q = mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * 5+:5];
	// Trace: core/cvfpu/src/fpnew_fma.sv:488:3
	wire [LOWER_SUM_WIDTH - 1:0] sum_lower;
	// Trace: core/cvfpu/src/fpnew_fma.sv:489:3
	wire [LZC_RESULT_WIDTH - 1:0] leading_zero_count;
	// Trace: core/cvfpu/src/fpnew_fma.sv:490:3
	wire signed [LZC_RESULT_WIDTH:0] leading_zero_count_sgn;
	// Trace: core/cvfpu/src/fpnew_fma.sv:491:3
	wire lzc_zeroes;
	// Trace: core/cvfpu/src/fpnew_fma.sv:493:3
	reg [SHIFT_AMOUNT_WIDTH - 1:0] norm_shamt;
	// Trace: core/cvfpu/src/fpnew_fma.sv:494:3
	reg signed [EXP_WIDTH - 1:0] normalized_exponent;
	// Trace: core/cvfpu/src/fpnew_fma.sv:496:3
	wire [(3 * PRECISION_BITS) + 4:0] sum_shifted;
	// Trace: core/cvfpu/src/fpnew_fma.sv:497:3
	reg [PRECISION_BITS:0] final_mantissa;
	// Trace: core/cvfpu/src/fpnew_fma.sv:498:3
	reg [(2 * PRECISION_BITS) + 2:0] sum_sticky_bits;
	// Trace: core/cvfpu/src/fpnew_fma.sv:499:3
	wire sticky_after_norm;
	// Trace: core/cvfpu/src/fpnew_fma.sv:501:3
	reg signed [EXP_WIDTH - 1:0] final_exponent;
	// Trace: core/cvfpu/src/fpnew_fma.sv:503:3
	assign sum_lower = sum_q[LOWER_SUM_WIDTH - 1:0];
	// Trace: core/cvfpu/src/fpnew_fma.sv:506:3
	lzc #(
		.WIDTH(LOWER_SUM_WIDTH),
		.MODE(1)
	) i_lzc(
		.in_i(sum_lower),
		.cnt_o(leading_zero_count),
		.empty_o(lzc_zeroes)
	);
	// Trace: core/cvfpu/src/fpnew_fma.sv:515:3
	assign leading_zero_count_sgn = $signed({1'b0, leading_zero_count});
	// Trace: core/cvfpu/src/fpnew_fma.sv:518:3
	always @(*) begin : norm_shift_amount
		if (_sv2v_0)
			;
		// Trace: core/cvfpu/src/fpnew_fma.sv:520:5
		if ((exponent_difference_q <= 0) || (effective_subtraction_q && (exponent_difference_q <= 2))) begin
			begin
				// Trace: core/cvfpu/src/fpnew_fma.sv:522:7
				if ((((exponent_product_q - leading_zero_count_sgn) + 1) >= 0) && !lzc_zeroes) begin
					// Trace: core/cvfpu/src/fpnew_fma.sv:524:9
					norm_shamt = (PRECISION_BITS + 2) + leading_zero_count;
					// Trace: core/cvfpu/src/fpnew_fma.sv:525:9
					normalized_exponent = (exponent_product_q - leading_zero_count_sgn) + 1;
				end
				else begin
					// Trace: core/cvfpu/src/fpnew_fma.sv:529:9
					norm_shamt = $unsigned(($signed(PRECISION_BITS) + 2) + exponent_product_q);
					// Trace: core/cvfpu/src/fpnew_fma.sv:530:9
					normalized_exponent = 0;
				end
			end
		end
		else begin
			// Trace: core/cvfpu/src/fpnew_fma.sv:534:7
			norm_shamt = addend_shamt_q;
			// Trace: core/cvfpu/src/fpnew_fma.sv:535:7
			normalized_exponent = tentative_exponent_q;
		end
	end
	// Trace: core/cvfpu/src/fpnew_fma.sv:540:3
	assign sum_shifted = sum_q << norm_shamt;
	// Trace: core/cvfpu/src/fpnew_fma.sv:544:3
	always @(*) begin : small_norm
		if (_sv2v_0)
			;
		// Trace: core/cvfpu/src/fpnew_fma.sv:546:5
		{final_mantissa, sum_sticky_bits} = sum_shifted;
		// Trace: core/cvfpu/src/fpnew_fma.sv:547:5
		final_exponent = normalized_exponent;
		// Trace: core/cvfpu/src/fpnew_fma.sv:550:5
		if (sum_shifted[(3 * PRECISION_BITS) + 4]) begin
			// Trace: core/cvfpu/src/fpnew_fma.sv:551:7
			{final_mantissa, sum_sticky_bits} = sum_shifted >> 1;
			// Trace: core/cvfpu/src/fpnew_fma.sv:552:7
			final_exponent = normalized_exponent + 1;
		end
		else if (sum_shifted[(3 * PRECISION_BITS) + 3])
			;
		else if (normalized_exponent > 1) begin
			// Trace: core/cvfpu/src/fpnew_fma.sv:558:7
			{final_mantissa, sum_sticky_bits} = sum_shifted << 1;
			// Trace: core/cvfpu/src/fpnew_fma.sv:559:7
			final_exponent = normalized_exponent - 1;
		end
		else
			// Trace: core/cvfpu/src/fpnew_fma.sv:562:7
			final_exponent = 1'sb0;
	end
	// Trace: core/cvfpu/src/fpnew_fma.sv:567:3
	assign sticky_after_norm = |{sum_sticky_bits} | sticky_before_add_q;
	// Trace: core/cvfpu/src/fpnew_fma.sv:572:3
	wire pre_round_sign;
	// Trace: core/cvfpu/src/fpnew_fma.sv:573:3
	wire [EXP_BITS - 1:0] pre_round_exponent;
	// Trace: core/cvfpu/src/fpnew_fma.sv:574:3
	wire [MAN_BITS - 1:0] pre_round_mantissa;
	// Trace: core/cvfpu/src/fpnew_fma.sv:575:3
	wire [(EXP_BITS + MAN_BITS) - 1:0] pre_round_abs;
	// Trace: core/cvfpu/src/fpnew_fma.sv:576:3
	wire [1:0] round_sticky_bits;
	// Trace: core/cvfpu/src/fpnew_fma.sv:578:3
	wire of_before_round;
	wire of_after_round;
	// Trace: core/cvfpu/src/fpnew_fma.sv:579:3
	wire uf_before_round;
	wire uf_after_round;
	// Trace: core/cvfpu/src/fpnew_fma.sv:580:3
	wire result_zero;
	// Trace: core/cvfpu/src/fpnew_fma.sv:582:3
	wire rounded_sign;
	// Trace: core/cvfpu/src/fpnew_fma.sv:583:3
	wire [(EXP_BITS + MAN_BITS) - 1:0] rounded_abs;
	// Trace: core/cvfpu/src/fpnew_fma.sv:586:3
	assign of_before_round = final_exponent >= ((2 ** EXP_BITS) - 1);
	// Trace: core/cvfpu/src/fpnew_fma.sv:587:3
	assign uf_before_round = final_exponent == 0;
	// Trace: core/cvfpu/src/fpnew_fma.sv:590:3
	assign pre_round_sign = final_sign_q;
	// Trace: core/cvfpu/src/fpnew_fma.sv:591:3
	assign pre_round_exponent = (of_before_round ? (2 ** EXP_BITS) - 2 : $unsigned(final_exponent[EXP_BITS - 1:0]));
	// Trace: core/cvfpu/src/fpnew_fma.sv:592:3
	assign pre_round_mantissa = (of_before_round ? {MAN_BITS {1'sb1}} : final_mantissa[MAN_BITS:1]);
	// Trace: core/cvfpu/src/fpnew_fma.sv:593:3
	assign pre_round_abs = {pre_round_exponent, pre_round_mantissa};
	// Trace: core/cvfpu/src/fpnew_fma.sv:596:3
	assign round_sticky_bits = (of_before_round ? 2'b11 : {final_mantissa[0], sticky_after_norm});
	// Trace: core/cvfpu/src/fpnew_fma.sv:599:3
	fpnew_rounding #(.AbsWidth(EXP_BITS + MAN_BITS)) i_fpnew_rounding(
		.abs_value_i(pre_round_abs),
		.sign_i(pre_round_sign),
		.round_sticky_bits_i(round_sticky_bits),
		.rnd_mode_i(rnd_mode_q),
		.effective_subtraction_i(effective_subtraction_q),
		.abs_rounded_o(rounded_abs),
		.sign_o(rounded_sign),
		.exact_zero_o(result_zero)
	);
	// Trace: core/cvfpu/src/fpnew_fma.sv:613:3
	assign uf_after_round = rounded_abs[(EXP_BITS + MAN_BITS) - 1:MAN_BITS] == {(((EXP_BITS + MAN_BITS) - 1) >= MAN_BITS ? (((EXP_BITS + MAN_BITS) - 1) - MAN_BITS) + 1 : (MAN_BITS - ((EXP_BITS + MAN_BITS) - 1)) + 1) * 1 {1'sb0}};
	// Trace: core/cvfpu/src/fpnew_fma.sv:614:3
	assign of_after_round = rounded_abs[(EXP_BITS + MAN_BITS) - 1:MAN_BITS] == {(((EXP_BITS + MAN_BITS) - 1) >= MAN_BITS ? (((EXP_BITS + MAN_BITS) - 1) - MAN_BITS) + 1 : (MAN_BITS - ((EXP_BITS + MAN_BITS) - 1)) + 1) * 1 {1'sb1}};
	// Trace: core/cvfpu/src/fpnew_fma.sv:619:3
	wire [WIDTH - 1:0] regular_result;
	// Trace: core/cvfpu/src/fpnew_fma.sv:620:3
	wire [4:0] regular_status;
	// Trace: core/cvfpu/src/fpnew_fma.sv:623:3
	assign regular_result = {rounded_sign, rounded_abs};
	// Trace: core/cvfpu/src/fpnew_fma.sv:624:3
	assign regular_status[4] = 1'b0;
	// Trace: core/cvfpu/src/fpnew_fma.sv:625:3
	assign regular_status[3] = 1'b0;
	// Trace: core/cvfpu/src/fpnew_fma.sv:626:3
	assign regular_status[2] = of_before_round | of_after_round;
	// Trace: core/cvfpu/src/fpnew_fma.sv:627:3
	assign regular_status[1] = uf_after_round & regular_status[0];
	// Trace: core/cvfpu/src/fpnew_fma.sv:628:3
	assign regular_status[0] = (|round_sticky_bits | of_before_round) | of_after_round;
	// Trace: core/cvfpu/src/fpnew_fma.sv:631:3
	wire [((1 + EXP_BITS) + MAN_BITS) - 1:0] result_d;
	// Trace: core/cvfpu/src/fpnew_fma.sv:632:3
	wire [4:0] status_d;
	// Trace: core/cvfpu/src/fpnew_fma.sv:635:3
	assign result_d = (result_is_special_q ? special_result_q : regular_result);
	// Trace: core/cvfpu/src/fpnew_fma.sv:636:3
	assign status_d = (result_is_special_q ? special_status_q : regular_status);
	// Trace: core/cvfpu/src/fpnew_fma.sv:642:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * ((1 + EXP_BITS) + MAN_BITS)) + ((NUM_OUT_REGS * ((1 + EXP_BITS) + MAN_BITS)) - 1) : ((NUM_OUT_REGS + 1) * ((1 + EXP_BITS) + MAN_BITS)) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * ((1 + EXP_BITS) + MAN_BITS) : 0)] out_pipe_result_q;
	// Trace: core/cvfpu/src/fpnew_fma.sv:643:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * 5) + ((NUM_OUT_REGS * 5) - 1) : ((NUM_OUT_REGS + 1) * 5) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * 5 : 0)] out_pipe_status_q;
	// Trace: core/cvfpu/src/fpnew_fma.sv:644:3
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + ((NUM_OUT_REGS * TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) - 1) : ((NUM_OUT_REGS + 1) * TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] : 0)] out_pipe_tag_q;
	// Trace: core/cvfpu/src/fpnew_fma.sv:645:3
	reg [0:NUM_OUT_REGS] out_pipe_mask_q;
	// Trace: core/cvfpu/src/fpnew_fma.sv:646:3
	reg [0:NUM_OUT_REGS] out_pipe_aux_q;
	// Trace: core/cvfpu/src/fpnew_fma.sv:647:3
	reg [0:NUM_OUT_REGS] out_pipe_valid_q;
	// Trace: core/cvfpu/src/fpnew_fma.sv:649:3
	wire [0:NUM_OUT_REGS] out_pipe_ready;
	// Trace: core/cvfpu/src/fpnew_fma.sv:652:3
	wire [((1 + EXP_BITS) + MAN_BITS) * 1:1] sv2v_tmp_4232B;
	assign sv2v_tmp_4232B = result_d;
	always @(*) out_pipe_result_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] = sv2v_tmp_4232B;
	// Trace: core/cvfpu/src/fpnew_fma.sv:653:3
	wire [5:1] sv2v_tmp_07934;
	assign sv2v_tmp_07934 = status_d;
	always @(*) out_pipe_status_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * 5+:5] = sv2v_tmp_07934;
	// Trace: core/cvfpu/src/fpnew_fma.sv:654:3
	wire [TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] * 1:1] sv2v_tmp_7C8F0;
	assign sv2v_tmp_7C8F0 = mid_pipe_tag_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]+:TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]];
	always @(*) out_pipe_tag_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]+:TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]] = sv2v_tmp_7C8F0;
	// Trace: core/cvfpu/src/fpnew_fma.sv:655:3
	wire [1:1] sv2v_tmp_D6E81;
	assign sv2v_tmp_D6E81 = mid_pipe_mask_q[NUM_MID_REGS];
	always @(*) out_pipe_mask_q[0] = sv2v_tmp_D6E81;
	// Trace: core/cvfpu/src/fpnew_fma.sv:656:3
	wire [1:1] sv2v_tmp_F4A83;
	assign sv2v_tmp_F4A83 = mid_pipe_aux_q[NUM_MID_REGS];
	always @(*) out_pipe_aux_q[0] = sv2v_tmp_F4A83;
	// Trace: core/cvfpu/src/fpnew_fma.sv:657:3
	wire [1:1] sv2v_tmp_E45E7;
	assign sv2v_tmp_E45E7 = mid_pipe_valid_q[NUM_MID_REGS];
	always @(*) out_pipe_valid_q[0] = sv2v_tmp_E45E7;
	// Trace: core/cvfpu/src/fpnew_fma.sv:659:3
	assign mid_pipe_ready[NUM_MID_REGS] = out_pipe_ready[0];
	// Trace: core/cvfpu/src/fpnew_fma.sv:661:3
	genvar _gv_i_68;
	generate
		for (_gv_i_68 = 0; _gv_i_68 < NUM_OUT_REGS; _gv_i_68 = _gv_i_68 + 1) begin : gen_output_pipeline
			localparam i = _gv_i_68;
			// Trace: core/cvfpu/src/fpnew_fma.sv:663:5
			wire reg_ena;
			// Trace: core/cvfpu/src/fpnew_fma.sv:667:5
			assign out_pipe_ready[i] = out_pipe_ready[i + 1] | ~out_pipe_valid_q[i + 1];
			// Trace: macro expansion of FFLARNC at core/cvfpu/src/fpnew_fma.sv:669:329
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFLARNC at core/cvfpu/src/fpnew_fma.sv:669:407
				if (!rst_ni)
					// Trace: macro expansion of FFLARNC at core/cvfpu/src/fpnew_fma.sv:669:485
					out_pipe_valid_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFLARNC at core/cvfpu/src/fpnew_fma.sv:669:637
					out_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (out_pipe_ready[i] ? out_pipe_valid_q[i] : out_pipe_valid_q[i + 1]));
			// Trace: core/cvfpu/src/fpnew_fma.sv:671:5
			assign reg_ena = out_pipe_ready[i] & out_pipe_valid_q[i];
			// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:673:67
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:673:164
				if (!rst_ni)
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:673:261
					out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:673:451
					out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] <= (reg_ena ? out_pipe_result_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] : out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS]);
			// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:674:67
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:674:164
				if (!rst_ni)
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:674:261
					out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:674:451
					out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= (reg_ena ? out_pipe_status_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * 5+:5] : out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5]);
			// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:675:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:675:174
				if (!rst_ni)
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:675:271
					out_pipe_tag_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]+:TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]] <= sv2v_cast_65D85(1'sb0);
				else
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:675:461
					out_pipe_tag_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]+:TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]] <= (reg_ena ? out_pipe_tag_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]+:TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]] : out_pipe_tag_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]+:TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]]);
			// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:676:67
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:676:164
				if (!rst_ni)
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:676:261
					out_pipe_mask_q[i + 1] <= 1'sb0;
				else
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:676:451
					out_pipe_mask_q[i + 1] <= (reg_ena ? out_pipe_mask_q[i] : out_pipe_mask_q[i + 1]);
			// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:677:77
			always @(posedge clk_i or negedge rst_ni)
				// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:677:174
				if (!rst_ni)
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:677:271
					out_pipe_aux_q[i + 1] <= 1'b0;
				else
					// Trace: macro expansion of FFL at core/cvfpu/src/fpnew_fma.sv:677:461
					out_pipe_aux_q[i + 1] <= (reg_ena ? out_pipe_aux_q[i] : out_pipe_aux_q[i + 1]);
		end
	endgenerate
	// Trace: core/cvfpu/src/fpnew_fma.sv:680:3
	assign out_pipe_ready[NUM_OUT_REGS] = out_ready_i;
	// Trace: core/cvfpu/src/fpnew_fma.sv:682:3
	assign result_o = out_pipe_result_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS];
	// Trace: core/cvfpu/src/fpnew_fma.sv:683:3
	assign status_o = out_pipe_status_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * 5+:5];
	// Trace: core/cvfpu/src/fpnew_fma.sv:684:3
	assign extension_bit_o = 1'b1;
	// Trace: core/cvfpu/src/fpnew_fma.sv:685:3
	assign tag_o = out_pipe_tag_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]+:TagType_TagType_TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]];
	// Trace: core/cvfpu/src/fpnew_fma.sv:686:3
	assign mask_o = out_pipe_mask_q[NUM_OUT_REGS];
	// Trace: core/cvfpu/src/fpnew_fma.sv:687:3
	assign aux_o = out_pipe_aux_q[NUM_OUT_REGS];
	// Trace: core/cvfpu/src/fpnew_fma.sv:688:3
	assign out_valid_o = out_pipe_valid_q[NUM_OUT_REGS];
	// Trace: core/cvfpu/src/fpnew_fma.sv:689:3
	assign busy_o = |{inp_pipe_valid_q, mid_pipe_valid_q, out_pipe_valid_q};
	initial _sv2v_0 = 0;
endmodule
