module hwpf_stride_wrapper_6E38E_28CF5 (
	clk_i,
	rst_ni,
	hwpf_stride_base_set_i,
	hwpf_stride_base_i,
	hwpf_stride_base_o,
	hwpf_stride_param_set_i,
	hwpf_stride_param_i,
	hwpf_stride_param_o,
	hwpf_stride_throttle_set_i,
	hwpf_stride_throttle_i,
	hwpf_stride_throttle_o,
	hwpf_stride_status_o,
	snoop_valid_i,
	snoop_abort_i,
	snoop_addr_offset_i,
	snoop_addr_tag_i,
	snoop_phys_indexed_i,
	hpdcache_req_sid_i,
	hpdcache_req_valid_o,
	hpdcache_req_ready_i,
	hpdcache_req_o,
	hpdcache_req_abort_o,
	hpdcache_req_tag_o,
	hpdcache_req_pma_o,
	hpdcache_rsp_valid_i,
	hpdcache_rsp_i
);
	// removed localparam type hpdcache_req_be_t_hpdcache_req_be_t_HPDcacheCfg_type
	parameter [1349:0] hpdcache_req_be_t_hpdcache_req_be_t_HPDcacheCfg = 0;
	// removed localparam type hpdcache_req_data_t_hpdcache_req_data_t_HPDcacheCfg_type
	parameter [1349:0] hpdcache_req_data_t_hpdcache_req_data_t_HPDcacheCfg = 0;
	// removed localparam type hpdcache_req_offset_t_hpdcache_req_offset_t_HPDcacheCfg_type
	parameter [1349:0] hpdcache_req_offset_t_hpdcache_req_offset_t_HPDcacheCfg = 0;
	// removed localparam type hpdcache_req_sid_t_hpdcache_req_sid_t_HPDcacheCfg_type
	parameter [1349:0] hpdcache_req_sid_t_hpdcache_req_sid_t_HPDcacheCfg = 0;
	// removed localparam type hpdcache_req_t_hpdcache_req_t_HPDcacheCfg_type
	parameter [1349:0] hpdcache_req_t_hpdcache_req_t_HPDcacheCfg = 0;
	// removed localparam type hpdcache_req_tid_t_hpdcache_req_tid_t_HPDcacheCfg_type
	parameter [1349:0] hpdcache_req_tid_t_hpdcache_req_tid_t_HPDcacheCfg = 0;
	// removed localparam type hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg_type
	parameter [1349:0] hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg = 0;
	// removed localparam type hpdcache_tag_t_hpdcache_tag_t_HPDcacheCfg_type
	parameter [1349:0] hpdcache_tag_t_hpdcache_tag_t_HPDcacheCfg = 0;
	reg _sv2v_0;
	// removed import hwpf_stride_pkg::*;
	// removed import hpdcache_pkg::*;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:34:15
	// removed localparam type hpdcache_pkg_hpdcache_victim_sel_policy_t
	// removed localparam type hpdcache_pkg_hpdcache_user_cfg_t
	// removed localparam type hpdcache_pkg_hpdcache_cfg_t
	parameter [1349:0] HPDcacheCfg = 1'sb0;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:35:15
	parameter [31:0] NUM_HW_PREFETCH = 4;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:36:15
	parameter [31:0] NUM_SNOOP_PORTS = 1;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:40:20
	// removed localparam type hpdcache_tag_t
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:41:20
	// removed localparam type hpdcache_req_offset_t
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:42:20
	// removed localparam type hpdcache_req_data_t
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:43:20
	// removed localparam type hpdcache_req_be_t
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:44:20
	// removed localparam type hpdcache_req_sid_t
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:45:20
	// removed localparam type hpdcache_req_tid_t
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:46:20
	// removed localparam type hpdcache_req_t
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:47:20
	// removed localparam type hpdcache_rsp_t
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:55:5
	input wire clk_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:56:5
	input wire rst_ni;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:60:5
	input wire [NUM_HW_PREFETCH - 1:0] hwpf_stride_base_set_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:61:5
	// removed localparam type hwpf_stride_pkg_hwpf_stride_base_t
	input wire [(NUM_HW_PREFETCH * 64) - 1:0] hwpf_stride_base_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:62:5
	output wire [(NUM_HW_PREFETCH * 64) - 1:0] hwpf_stride_base_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:64:5
	input wire [NUM_HW_PREFETCH - 1:0] hwpf_stride_param_set_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:65:5
	// removed localparam type hwpf_stride_pkg_hwpf_stride_param_t
	input wire [(NUM_HW_PREFETCH * 64) - 1:0] hwpf_stride_param_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:66:5
	output wire [(NUM_HW_PREFETCH * 64) - 1:0] hwpf_stride_param_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:68:5
	input wire [NUM_HW_PREFETCH - 1:0] hwpf_stride_throttle_set_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:69:5
	// removed localparam type hwpf_stride_pkg_hwpf_stride_throttle_t
	input wire [(NUM_HW_PREFETCH * 32) - 1:0] hwpf_stride_throttle_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:70:5
	output wire [(NUM_HW_PREFETCH * 32) - 1:0] hwpf_stride_throttle_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:72:5
	// removed localparam type hwpf_stride_pkg_hwpf_stride_status_t
	output wire [63:0] hwpf_stride_status_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:77:5
	input wire [NUM_SNOOP_PORTS - 1:0] snoop_valid_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:78:5
	input wire [NUM_SNOOP_PORTS - 1:0] snoop_abort_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:79:5
	input wire [(NUM_SNOOP_PORTS * hpdcache_req_offset_t_hpdcache_req_offset_t_HPDcacheCfg[287-:32]) - 1:0] snoop_addr_offset_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:80:5
	input wire [(NUM_SNOOP_PORTS * hpdcache_tag_t_hpdcache_tag_t_HPDcacheCfg[351-:32]) - 1:0] snoop_addr_tag_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:81:5
	input wire [NUM_SNOOP_PORTS - 1:0] snoop_phys_indexed_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:86:5
	input wire [hpdcache_req_sid_t_hpdcache_req_sid_t_HPDcacheCfg[1093-:32] - 1:0] hpdcache_req_sid_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:87:5
	output wire hpdcache_req_valid_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:88:5
	input wire hpdcache_req_ready_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:89:5
	output wire [((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1:0] hpdcache_req_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:90:5
	output wire hpdcache_req_abort_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:91:5
	output wire [hpdcache_tag_t_hpdcache_tag_t_HPDcacheCfg[351-:32] - 1:0] hpdcache_req_tag_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:92:5
	// removed localparam type hpdcache_pkg_hpdcache_pma_t
	output wire [1:0] hpdcache_req_pma_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:93:5
	input wire hpdcache_rsp_valid_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:94:5
	input wire [(((hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1157-:32] * hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1285-:32]) + hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32]) + hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32]) + 1:0] hpdcache_rsp_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:101:5
	// removed localparam type hpdcache_nline_t
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:102:5
	// removed localparam type hpdcache_set_t
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:107:5
	reg [NUM_SNOOP_PORTS - 1:0] snoop_valid_q;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:108:5
	reg [(NUM_SNOOP_PORTS * hpdcache_req_offset_t_hpdcache_req_offset_t_HPDcacheCfg[287-:32]) - 1:0] snoop_addr_offset_q;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:113:5
	wire [NUM_HW_PREFETCH - 1:0] hwpf_stride_enable;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:114:5
	wire [NUM_HW_PREFETCH - 1:0] hwpf_stride_free;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:115:5
	wire [NUM_HW_PREFETCH - 1:0] hwpf_stride_status_busy;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:116:5
	reg [3:0] hwpf_stride_status_free_idx;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:118:5
	wire [(NUM_HW_PREFETCH * HPDcacheCfg[383-:32]) - 1:0] hwpf_snoop_nline;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:119:5
	reg [NUM_HW_PREFETCH - 1:0] hwpf_snoop_match;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:121:5
	wire [NUM_HW_PREFETCH - 1:0] hwpf_stride_req_valid;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:122:5
	wire [NUM_HW_PREFETCH - 1:0] hwpf_stride_req_ready;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:123:5
	wire [((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? (NUM_HW_PREFETCH * (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 2)) - 1 : (NUM_HW_PREFETCH * (1 - (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1))) + (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 0)):((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? 0 : ((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1)] hwpf_stride_req;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:125:5
	wire [NUM_HW_PREFETCH - 1:0] hwpf_stride_arb_in_req_valid;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:126:5
	wire [NUM_HW_PREFETCH - 1:0] hwpf_stride_arb_in_req_ready;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:127:5
	wire [((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? (NUM_HW_PREFETCH * (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 2)) - 1 : (NUM_HW_PREFETCH * (1 - (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1))) + (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 0)):((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? 0 : ((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1)] hwpf_stride_arb_in_req;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:128:5
	wire [NUM_HW_PREFETCH - 1:0] hwpf_stride_arb_in_rsp_valid;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:129:5
	wire [(((((hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1157-:32] * hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1285-:32]) + hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32]) + hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32]) + 1) >= 0 ? (NUM_HW_PREFETCH * ((((hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1157-:32] * hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1285-:32]) + hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32]) + hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32]) + 2)) - 1 : (NUM_HW_PREFETCH * (1 - ((((hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1157-:32] * hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1285-:32]) + hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32]) + hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32]) + 1))) + ((((hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1157-:32] * hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1285-:32]) + hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32]) + hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32]) + 0)):(((((hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1157-:32] * hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1285-:32]) + hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32]) + hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32]) + 1) >= 0 ? 0 : (((hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1157-:32] * hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1285-:32]) + hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32]) + hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32]) + 1)] hwpf_stride_arb_in_rsp;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:135:5
	initial begin : initial_assertions
		// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:137:9
		begin : max_hwpf_stride_assert
			
		end
	end
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:145:5
	always @(*) begin : sv2v_autoblock_1
		reg [0:1] _sv2v_jump;
		_sv2v_jump = 2'b00;
		begin : hwpf_stride_priority_encoder
			if (_sv2v_0)
				;
			// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:146:9
			hwpf_stride_status_free_idx = 1'sb0;
			// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:147:9
			begin : sv2v_autoblock_2
				// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:147:14
				reg [31:0] i;
				// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:147:14
				begin : sv2v_autoblock_3
					reg [31:0] _sv2v_value_on_break;
					for (i = 0; i < NUM_HW_PREFETCH; i = i + 1)
						if (_sv2v_jump < 2'b10) begin
							_sv2v_jump = 2'b00;
							// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:148:13
							if (hwpf_stride_free[i]) begin
								// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:149:17
								hwpf_stride_status_free_idx = i;
								// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:150:17
								_sv2v_jump = 2'b10;
							end
							_sv2v_value_on_break = i;
						end
					if (!(_sv2v_jump < 2'b10))
						i = _sv2v_value_on_break;
					if (_sv2v_jump != 2'b11)
						_sv2v_jump = 2'b00;
				end
			end
		end
	end
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:156:5
	assign hwpf_stride_free = ~(hwpf_stride_enable | hwpf_stride_status_busy);
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:158:5
	assign hwpf_stride_status_o[63:32] = {{32 - NUM_HW_PREFETCH {1'b0}}, hwpf_stride_status_busy};
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:160:5
	assign hwpf_stride_status_o[31] = |hwpf_stride_free;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:162:5
	assign hwpf_stride_status_o[30:16] = {11'b00000000000, hwpf_stride_status_free_idx};
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:164:5
	assign hwpf_stride_status_o[15:0] = {{16 - NUM_HW_PREFETCH {1'b0}}, hwpf_stride_enable};
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:169:5
	genvar _gv_j_12;
	generate
		for (_gv_j_12 = 0; _gv_j_12 < NUM_SNOOP_PORTS; _gv_j_12 = _gv_j_12 + 1) begin : gen_hwpf_snoop
			localparam j = _gv_j_12;
			// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:170:9
			always @(posedge clk_i or negedge rst_ni) begin : snoop_ff
				// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:172:13
				if (!rst_ni) begin
					// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:173:17
					snoop_valid_q[j] <= 1'b0;
					// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:174:17
					snoop_addr_offset_q[j * hpdcache_req_offset_t_hpdcache_req_offset_t_HPDcacheCfg[287-:32]+:hpdcache_req_offset_t_hpdcache_req_offset_t_HPDcacheCfg[287-:32]] <= 1'sb0;
				end
				else
					// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:176:17
					if (snoop_phys_indexed_i[j]) begin
						// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:177:21
						snoop_valid_q[j] <= snoop_valid_i[j];
						// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:178:21
						snoop_addr_offset_q[j * hpdcache_req_offset_t_hpdcache_req_offset_t_HPDcacheCfg[287-:32]+:hpdcache_req_offset_t_hpdcache_req_offset_t_HPDcacheCfg[287-:32]] <= snoop_addr_offset_i[j * hpdcache_req_offset_t_hpdcache_req_offset_t_HPDcacheCfg[287-:32]+:hpdcache_req_offset_t_hpdcache_req_offset_t_HPDcacheCfg[287-:32]];
					end
			end
		end
	endgenerate
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:184:5
	genvar _gv_i_80;
	function automatic [hpdcache_req_tid_t_hpdcache_req_tid_t_HPDcacheCfg[1125-:32] - 1:0] sv2v_cast_3A03B;
		input reg [hpdcache_req_tid_t_hpdcache_req_tid_t_HPDcacheCfg[1125-:32] - 1:0] inp;
		sv2v_cast_3A03B = inp;
	endfunction
	generate
		for (_gv_i_80 = 0; _gv_i_80 < NUM_HW_PREFETCH; _gv_i_80 = _gv_i_80 + 1) begin : gen_hwpf_stride
			localparam i = _gv_i_80;
			// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:185:9
			assign hwpf_stride_enable[i] = hwpf_stride_base_o[i * 64];
			// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:189:9
			always @(*) begin : snoop_comb
				if (_sv2v_0)
					;
				// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:191:13
				hwpf_snoop_match[i] = 1'b0;
				// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:192:13
				begin : sv2v_autoblock_4
					// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:192:18
					reg signed [31:0] j;
					// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:192:18
					for (j = 0; j < NUM_SNOOP_PORTS; j = j + 1)
						begin : sv2v_autoblock_5
							// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:193:17
							reg snoop_valid;
							// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:194:17
							reg [hpdcache_req_offset_t_hpdcache_req_offset_t_HPDcacheCfg[287-:32] - 1:0] snoop_offset;
							// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:195:17
							reg [HPDcacheCfg[383-:32] - 1:0] snoop_nline;
							// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:197:17
							if (snoop_phys_indexed_i[j]) begin
								// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:198:21
								snoop_valid = snoop_valid_i[j];
								// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:199:21
								snoop_offset = snoop_addr_offset_i[j * hpdcache_req_offset_t_hpdcache_req_offset_t_HPDcacheCfg[287-:32]+:hpdcache_req_offset_t_hpdcache_req_offset_t_HPDcacheCfg[287-:32]];
							end
							else begin
								// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:201:21
								snoop_valid = snoop_valid_q[j];
								// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:202:21
								snoop_offset = snoop_addr_offset_q[j * hpdcache_req_offset_t_hpdcache_req_offset_t_HPDcacheCfg[287-:32]+:hpdcache_req_offset_t_hpdcache_req_offset_t_HPDcacheCfg[287-:32]];
							end
							// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:204:17
							snoop_nline = {snoop_addr_tag_i[j * hpdcache_tag_t_hpdcache_tag_t_HPDcacheCfg[351-:32]+:hpdcache_tag_t_hpdcache_tag_t_HPDcacheCfg[351-:32]], snoop_offset};
							// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:205:17
							hwpf_snoop_match[i] = hwpf_snoop_match[i] | ((snoop_valid && !snoop_abort_i[j]) && (hwpf_snoop_nline[i * HPDcacheCfg[383-:32]+:HPDcacheCfg[383-:32]] == snoop_nline));
						end
				end
			end
			// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:211:9
			hwpf_stride_04E73_7B29C #(
				.hpdcache_nline_t_HPDcacheCfg(HPDcacheCfg),
				.hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg(hpdcache_req_t_hpdcache_req_t_HPDcacheCfg),
				.hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg(hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg),
				.hpdcache_set_t_HPDcacheCfg(HPDcacheCfg),
				.hpdcache_tag_t_hpdcache_tag_t_hpdcache_tag_t_HPDcacheCfg(hpdcache_tag_t_hpdcache_tag_t_HPDcacheCfg),
				.HPDcacheCfg(HPDcacheCfg)
			) hwpf_stride_i(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.csr_base_set_i(hwpf_stride_base_set_i[i]),
				.csr_base_i(hwpf_stride_base_i[i * 64+:64]),
				.csr_param_set_i(hwpf_stride_param_set_i[i]),
				.csr_param_i(hwpf_stride_param_i[i * 64+:64]),
				.csr_throttle_set_i(hwpf_stride_throttle_set_i[i]),
				.csr_throttle_i(hwpf_stride_throttle_i[i * 32+:32]),
				.csr_base_o(hwpf_stride_base_o[i * 64+:64]),
				.csr_param_o(hwpf_stride_param_o[i * 64+:64]),
				.csr_throttle_o(hwpf_stride_throttle_o[i * 32+:32]),
				.busy_o(hwpf_stride_status_busy[i]),
				.snoop_nline_o(hwpf_snoop_nline[i * HPDcacheCfg[383-:32]+:HPDcacheCfg[383-:32]]),
				.snoop_match_i(hwpf_snoop_match[i]),
				.hpdcache_req_valid_o(hwpf_stride_req_valid[i]),
				.hpdcache_req_ready_i(hwpf_stride_req_ready[i]),
				.hpdcache_req_o(hwpf_stride_req[((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? 0 : ((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) + (i * ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? ((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 2 : 1 - (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1)))+:((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? ((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 2 : 1 - (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1))]),
				.hpdcache_rsp_valid_i(hwpf_stride_arb_in_rsp_valid[i]),
				.hpdcache_rsp_i(hwpf_stride_arb_in_rsp[(((((hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1157-:32] * hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1285-:32]) + hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32]) + hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32]) + 1) >= 0 ? 0 : (((hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1157-:32] * hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1285-:32]) + hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32]) + hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32]) + 1) + (i * (((((hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1157-:32] * hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1285-:32]) + hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32]) + hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32]) + 1) >= 0 ? (((hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1157-:32] * hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1285-:32]) + hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32]) + hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32]) + 2 : 1 - ((((hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1157-:32] * hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1285-:32]) + hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32]) + hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32]) + 1)))+:(((((hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1157-:32] * hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1285-:32]) + hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32]) + hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32]) + 1) >= 0 ? (((hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1157-:32] * hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1285-:32]) + hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32]) + hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32]) + 2 : 1 - ((((hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1157-:32] * hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1285-:32]) + hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32]) + hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32]) + 1))])
			);
			// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:245:9
			assign hwpf_stride_req_ready[i] = hwpf_stride_arb_in_req_ready[i];
			assign hwpf_stride_arb_in_req_valid[i] = hwpf_stride_req_valid[i];
			assign hwpf_stride_arb_in_req[((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? (i * ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? ((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 2 : 1 - (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1))) + ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) : (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) - (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))))) : (((i * ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? ((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 2 : 1 - (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1))) + ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) : (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) - (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))))) + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))) >= ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))))) ? ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))) - ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))))) + 1 : (((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))))) - (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))))) + 1)) - 1)-:((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))) >= ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))))) ? ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))) - ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))))) + 1 : (((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))))) - (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))))) + 1)] = hwpf_stride_req[((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? (i * ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? ((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 2 : 1 - (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1))) + ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) : (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) - (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))))) : (((i * ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? ((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 2 : 1 - (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1))) + ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) : (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) - (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))))) + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))) >= ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))))) ? ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))) - ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))))) + 1 : (((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))))) - (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))))) + 1)) - 1)-:((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))) >= ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))))) ? ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))) - ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))))) + 1 : (((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))))) - (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))))) + 1)];
			assign hwpf_stride_arb_in_req[((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? (i * ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? ((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 2 : 1 - (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1))) + ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) : (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) - ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))) : (((i * ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? ((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 2 : 1 - (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1))) + ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) : (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) - ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))))) + (((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) >= (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) ? (((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) - (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))))) + 1 : ((4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) - ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))) + 1)) - 1)-:(((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) >= (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) ? (((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) - (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))))) + 1 : ((4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) - ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))) + 1)] = hwpf_stride_req[((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? (i * ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? ((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 2 : 1 - (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1))) + ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) : (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) - ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))) : (((i * ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? ((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 2 : 1 - (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1))) + ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) : (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) - ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))))) + (((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) >= (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) ? (((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) - (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))))) + 1 : ((4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) - ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))) + 1)) - 1)-:(((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) >= (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) ? (((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) - (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))))) + 1 : ((4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) - ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))) + 1)];
			assign hwpf_stride_arb_in_req[((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? (i * ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? ((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 2 : 1 - (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1))) + ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? 4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) : (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) - (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) : (((i * ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? ((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 2 : 1 - (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1))) + ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? 4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) : (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) - (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))) + ((4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) >= ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) ? ((4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) - ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) + 1 : (((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) - (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) + 1)) - 1)-:((4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) >= ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) ? ((4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) - ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) + 1 : (((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) - (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) + 1)] = hwpf_stride_req[((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? (i * ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? ((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 2 : 1 - (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1))) + ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? 4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) : (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) - (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) : (((i * ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? ((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 2 : 1 - (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1))) + ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? 4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) : (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) - (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))) + ((4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) >= ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) ? ((4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) - ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) + 1 : (((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) - (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) + 1)) - 1)-:((4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) >= ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) ? ((4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) - ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) + 1 : (((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) - (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) + 1)];
			assign hwpf_stride_arb_in_req[((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? (i * ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? ((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 2 : 1 - (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1))) + ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) : (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) - ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) : (((i * ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? ((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 2 : 1 - (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1))) + ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) : (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) - ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) + (((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) >= (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))) ? (((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) - (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) + 1 : ((3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))) - ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) + 1)) - 1)-:(((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) >= (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))) ? (((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) - (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) + 1 : ((3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))) - ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) + 1)] = hwpf_stride_req[((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? (i * ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? ((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 2 : 1 - (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1))) + ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) : (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) - ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) : (((i * ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? ((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 2 : 1 - (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1))) + ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) : (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) - ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) + (((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) >= (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))) ? (((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) - (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) + 1 : ((3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))) - ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) + 1)) - 1)-:(((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) >= (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))) ? (((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) - (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) + 1 : ((3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))) - ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) + 1)];
			assign hwpf_stride_arb_in_req[((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? (i * ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? ((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 2 : 1 - (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1))) + ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? 3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))) : (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) - (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) : (((i * ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? ((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 2 : 1 - (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1))) + ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? 3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))) : (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) - (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) + ((3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) >= (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) ? ((3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) - (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))) + 1 : ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) - (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) + 1)) - 1)-:((3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) >= (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) ? ((3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) - (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))) + 1 : ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) - (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) + 1)] = hwpf_stride_req[((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? (i * ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? ((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 2 : 1 - (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1))) + ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? 3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))) : (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) - (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) : (((i * ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? ((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 2 : 1 - (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1))) + ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? 3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))) : (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) - (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) + ((3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) >= (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) ? ((3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) - (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))) + 1 : ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) - (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) + 1)) - 1)-:((3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) >= (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) ? ((3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) - (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))) + 1 : ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) - (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) + 1)];
			assign hwpf_stride_arb_in_req[((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? (i * ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? ((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 2 : 1 - (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1))) + ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))) : (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) - (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) : (((i * ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? ((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 2 : 1 - (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1))) + ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))) : (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) - (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))) >= (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))) ? ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))) - (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) + 1 : ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))) - (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) + 1)) - 1)-:((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))) >= (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))) ? ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))) - (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) + 1 : ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))) - (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) + 1)] = hpdcache_req_sid_i;
			assign hwpf_stride_arb_in_req[((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? (i * ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? ((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 2 : 1 - (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1))) + ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)) : (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) - (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))) : (((i * ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? ((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 2 : 1 - (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1))) + ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)) : (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) - (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))) >= (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)) ? ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))) - (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))) + 1 : ((2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)) - (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))) + 1)) - 1)-:((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))) >= (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)) ? ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))) - (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))) + 1 : ((2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)) - (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))) + 1)] = sv2v_cast_3A03B(i);
			assign hwpf_stride_arb_in_req[(i * ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? ((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 2 : 1 - (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1))) + ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? 2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1) : (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) - (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))] = hwpf_stride_req[(i * ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? ((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 2 : 1 - (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1))) + ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? 2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1) : (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) - (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))];
			assign hwpf_stride_arb_in_req[(i * ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? ((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 2 : 1 - (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1))) + ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? 1 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1) : (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) - (1 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))] = hwpf_stride_req[(i * ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? ((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 2 : 1 - (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1))) + ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? 1 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1) : (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) - (1 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))];
			assign hwpf_stride_arb_in_req[((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? (i * ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? ((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 2 : 1 - (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1))) + ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1 : (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) - (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)) : (((i * ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? ((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 2 : 1 - (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1))) + ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1 : (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) - (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))) + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1) >= 2 ? hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 0 : 3 - (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))) - 1)-:((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1) >= 2 ? hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 0 : 3 - (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))] = 1'sb0;
			assign hwpf_stride_arb_in_req[((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? (i * ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? ((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 2 : 1 - (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1))) + ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? 1 : ((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 0) : ((i * ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? ((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 2 : 1 - (((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1))) + ((((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1) >= 0 ? 1 : ((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 0)) + 1)-:2] = 1'sb0;
		end
	endgenerate
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:263:5
	hwpf_stride_arb_47A89_10D5A #(
		.hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg(hpdcache_req_t_hpdcache_req_t_HPDcacheCfg),
		.hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg(hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg),
		.NUM_HW_PREFETCH(NUM_HW_PREFETCH)
	) hwpf_stride_arb_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.hwpf_stride_req_valid_i(hwpf_stride_arb_in_req_valid),
		.hwpf_stride_req_ready_o(hwpf_stride_arb_in_req_ready),
		.hwpf_stride_req_i(hwpf_stride_arb_in_req),
		.hwpf_stride_rsp_valid_o(hwpf_stride_arb_in_rsp_valid),
		.hwpf_stride_rsp_o(hwpf_stride_arb_in_rsp),
		.hpdcache_req_valid_o(hpdcache_req_valid_o),
		.hpdcache_req_ready_i(hpdcache_req_ready_i),
		.hpdcache_req_o(hpdcache_req_o),
		.hpdcache_rsp_valid_i(hpdcache_rsp_valid_i),
		.hpdcache_rsp_i(hpdcache_rsp_i)
	);
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hwpf_stride/hwpf_stride_wrapper.sv:286:5
	assign hpdcache_req_abort_o = 1'b0;
	assign hpdcache_req_tag_o = 1'sb0;
	assign hpdcache_req_pma_o = 1'sb0;
	initial _sv2v_0 = 0;
endmodule
