module hpdcache_mem_to_axi_write_A24E0_6C8C1 (
	req_ready_o,
	req_valid_i,
	req_i,
	req_data_ready_o,
	req_data_valid_i,
	req_data_i,
	resp_ready_i,
	resp_valid_o,
	resp_o,
	axi_aw_valid_o,
	axi_aw_o,
	axi_aw_ready_i,
	axi_w_valid_o,
	axi_w_o,
	axi_w_ready_i,
	axi_b_valid_i,
	axi_b_i,
	axi_b_ready_o
);
	// removed localparam type aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_AddrWidth_type
	// removed localparam type aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_IdWidth_type
	// removed localparam type aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth_type
	parameter signed [31:0] aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_AddrWidth = 0;
	parameter signed [31:0] aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_IdWidth = 0;
	parameter signed [31:0] aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth = 0;
	// removed localparam type b_chan_t_axi_b_chan_t_axi_b_chan_t_CVA6Cfg_type
	// removed localparam type b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules_type
	parameter [17102:0] b_chan_t_axi_b_chan_t_axi_b_chan_t_CVA6Cfg = 0;
	parameter signed [31:0] b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules = 0;
	// removed localparam type hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg_type
	parameter [1349:0] hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg = 0;
	// removed localparam type hpdcache_mem_req_w_t_hpdcache_mem_req_w_t_HPDcacheCfg_type
	parameter [1349:0] hpdcache_mem_req_w_t_hpdcache_mem_req_w_t_HPDcacheCfg = 0;
	// removed localparam type hpdcache_mem_resp_w_t_hpdcache_mem_resp_w_t_HPDcacheCfg_type
	parameter [1349:0] hpdcache_mem_resp_w_t_hpdcache_mem_resp_w_t_HPDcacheCfg = 0;
	// removed localparam type w_chan_t_axi_w_chan_t_axi_w_chan_t_axi_w_chan_t_ariane_axi_DataWidth_type
	// removed localparam type w_chan_t_axi_w_chan_t_axi_w_chan_t_axi_w_chan_t_ariane_axi_StrbWidth_type
	// removed localparam type w_chan_t_axi_w_chan_t_axi_w_chan_t_axi_w_chan_t_ariane_axi_UserWidth_type
	parameter signed [31:0] w_chan_t_axi_w_chan_t_axi_w_chan_t_axi_w_chan_t_ariane_axi_DataWidth = 0;
	parameter signed [31:0] w_chan_t_axi_w_chan_t_axi_w_chan_t_axi_w_chan_t_ariane_axi_StrbWidth = 0;
	parameter signed [31:0] w_chan_t_axi_w_chan_t_axi_w_chan_t_axi_w_chan_t_ariane_axi_UserWidth = 0;
	reg _sv2v_0;
	// removed import hpdcache_pkg::*;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_write.sv:29:20
	// removed localparam type hpdcache_mem_req_t
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_write.sv:30:20
	// removed localparam type hpdcache_mem_req_w_t
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_write.sv:31:20
	// removed localparam type hpdcache_mem_resp_w_t
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_write.sv:32:20
	// removed localparam type aw_chan_t
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_write.sv:33:20
	// removed localparam type w_chan_t
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_write.sv:34:20
	// removed localparam type b_chan_t
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_write.sv:37:5
	output wire req_ready_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_write.sv:38:5
	input wire req_valid_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_write.sv:39:5
	input wire [((hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[639-:32] + 11) + hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[607-:32]) + 6:0] req_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_write.sv:41:5
	output wire req_data_ready_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_write.sv:42:5
	input wire req_data_valid_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_write.sv:43:5
	input wire [(hpdcache_mem_req_w_t_hpdcache_mem_req_w_t_HPDcacheCfg[575-:32] + (hpdcache_mem_req_w_t_hpdcache_mem_req_w_t_HPDcacheCfg[575-:32] / 8)) + 0:0] req_data_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_write.sv:45:5
	input wire resp_ready_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_write.sv:46:5
	output wire resp_valid_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_write.sv:47:5
	output wire [(3 + hpdcache_mem_resp_w_t_hpdcache_mem_resp_w_t_HPDcacheCfg[607-:32]) - 1:0] resp_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_write.sv:49:5
	output wire axi_aw_valid_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_write.sv:50:5
	output wire [(((aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_IdWidth + aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_AddrWidth) + 35) + aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth) - 1:0] axi_aw_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_write.sv:51:5
	input wire axi_aw_ready_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_write.sv:53:5
	output wire axi_w_valid_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_write.sv:54:5
	output wire [(((w_chan_t_axi_w_chan_t_axi_w_chan_t_axi_w_chan_t_ariane_axi_DataWidth + w_chan_t_axi_w_chan_t_axi_w_chan_t_axi_w_chan_t_ariane_axi_StrbWidth) + 1) + w_chan_t_axi_w_chan_t_axi_w_chan_t_axi_w_chan_t_ariane_axi_UserWidth) - 1:0] axi_w_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_write.sv:55:5
	input wire axi_w_ready_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_write.sv:57:5
	input wire axi_b_valid_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_write.sv:58:5
	input wire [((b_chan_t_axi_b_chan_t_axi_b_chan_t_CVA6Cfg[9119 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9119 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9119 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9119 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 2) + b_chan_t_axi_b_chan_t_axi_b_chan_t_CVA6Cfg[9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) - 1:0] axi_b_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_write.sv:59:5
	output wire axi_b_ready_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_write.sv:62:5
	reg lock;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_write.sv:63:5
	// removed localparam type axi_pkg_atop_t
	reg [5:0] atop;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_write.sv:64:5
	// removed localparam type axi_pkg_cache_t
	wire [3:0] cache;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_write.sv:65:5
	// removed localparam type hpdcache_pkg_hpdcache_mem_error_e
	reg [1:0] resp;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_write.sv:67:5
	localparam axi_pkg_ATOP_ADD = 3'b000;
	localparam axi_pkg_ATOP_ATOMICLOAD = 2'b10;
	localparam axi_pkg_ATOP_ATOMICSWAP = 6'b110000;
	localparam axi_pkg_ATOP_CLR = 3'b001;
	localparam axi_pkg_ATOP_EOR = 3'b010;
	localparam axi_pkg_ATOP_LITTLE_END = 1'b0;
	localparam axi_pkg_ATOP_SET = 3'b011;
	localparam axi_pkg_ATOP_SMAX = 3'b100;
	localparam axi_pkg_ATOP_SMIN = 3'b101;
	localparam axi_pkg_ATOP_UMAX = 3'b110;
	localparam axi_pkg_ATOP_UMIN = 3'b111;
	// removed localparam type hpdcache_pkg_hpdcache_mem_command_e
	// removed localparam type hpdcache_pkg_hpdcache_mem_atomic_e
	always @(*) begin : atop_comb
		if (_sv2v_0)
			;
		// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_write.sv:69:9
		lock = 1'b0;
		// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_write.sv:70:9
		atop = 1'sb0;
		// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_write.sv:71:9
		case (req_i[6-:2])
			2'b10:
				// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_write.sv:73:17
				case (req_i[4-:4])
					4'b1101:
						// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_write.sv:74:47
						lock = 1'b1;
					4'b0000:
						// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_write.sv:75:47
						atop = {axi_pkg_ATOP_ATOMICLOAD, axi_pkg_ATOP_LITTLE_END, axi_pkg_ATOP_ADD};
					4'b0001:
						// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_write.sv:78:47
						atop = {axi_pkg_ATOP_ATOMICLOAD, axi_pkg_ATOP_LITTLE_END, axi_pkg_ATOP_CLR};
					4'b0010:
						// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_write.sv:81:47
						atop = {axi_pkg_ATOP_ATOMICLOAD, axi_pkg_ATOP_LITTLE_END, axi_pkg_ATOP_SET};
					4'b0011:
						// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_write.sv:84:47
						atop = {axi_pkg_ATOP_ATOMICLOAD, axi_pkg_ATOP_LITTLE_END, axi_pkg_ATOP_EOR};
					4'b0100:
						// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_write.sv:87:47
						atop = {axi_pkg_ATOP_ATOMICLOAD, axi_pkg_ATOP_LITTLE_END, axi_pkg_ATOP_SMAX};
					4'b0101:
						// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_write.sv:90:47
						atop = {axi_pkg_ATOP_ATOMICLOAD, axi_pkg_ATOP_LITTLE_END, axi_pkg_ATOP_SMIN};
					4'b0110:
						// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_write.sv:93:47
						atop = {axi_pkg_ATOP_ATOMICLOAD, axi_pkg_ATOP_LITTLE_END, axi_pkg_ATOP_UMAX};
					4'b0111:
						// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_write.sv:96:47
						atop = {axi_pkg_ATOP_ATOMICLOAD, axi_pkg_ATOP_LITTLE_END, axi_pkg_ATOP_UMIN};
					4'b1000:
						// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_write.sv:99:47
						atop = axi_pkg_ATOP_ATOMICSWAP;
				endcase
		endcase
	end
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_write.sv:105:5
	localparam axi_pkg_CACHE_BUFFERABLE = 4'b0001;
	localparam axi_pkg_CACHE_MODIFIABLE = 4'b0010;
	localparam axi_pkg_CACHE_RD_ALLOC = 4'b0100;
	localparam axi_pkg_CACHE_WR_ALLOC = 4'b1000;
	assign cache = (req_i[0] && !lock ? ((axi_pkg_CACHE_BUFFERABLE | axi_pkg_CACHE_MODIFIABLE) | axi_pkg_CACHE_RD_ALLOC) | axi_pkg_CACHE_WR_ALLOC : {4 {1'sb0}});
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_write.sv:111:5
	localparam axi_pkg_RESP_DECERR = 2'b11;
	localparam axi_pkg_RESP_SLVERR = 2'b10;
	always @(*) begin : resp_decode_comb
		if (_sv2v_0)
			;
		// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_write.sv:113:9
		case (axi_b_i[b_chan_t_axi_b_chan_t_axi_b_chan_t_CVA6Cfg[9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 1-:((b_chan_t_axi_b_chan_t_axi_b_chan_t_CVA6Cfg[9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 1) >= (b_chan_t_axi_b_chan_t_axi_b_chan_t_CVA6Cfg[9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0) ? ((b_chan_t_axi_b_chan_t_axi_b_chan_t_CVA6Cfg[9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 1) - (b_chan_t_axi_b_chan_t_axi_b_chan_t_CVA6Cfg[9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0)) + 1 : ((b_chan_t_axi_b_chan_t_axi_b_chan_t_CVA6Cfg[9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0) - (b_chan_t_axi_b_chan_t_axi_b_chan_t_CVA6Cfg[9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 1)) + 1)])
			axi_pkg_RESP_SLVERR, axi_pkg_RESP_DECERR:
				// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_write.sv:115:35
				resp = 2'b01;
			default:
				// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_write.sv:116:35
				resp = 2'b00;
		endcase
	end
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_write.sv:120:5
	assign req_ready_o = axi_aw_ready_i;
	assign axi_aw_valid_o = req_valid_i;
	assign axi_aw_o[aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_IdWidth + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_AddrWidth + (29 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 5)))-:((aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_IdWidth + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_AddrWidth + (29 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 5)))) >= (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_AddrWidth + (35 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 0))) ? ((aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_IdWidth + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_AddrWidth + (29 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 5)))) - (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_AddrWidth + (35 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 0)))) + 1 : ((aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_AddrWidth + (35 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 0))) - (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_IdWidth + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_AddrWidth + (29 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 5))))) + 1)] = req_i[hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[607-:32] + 6-:((hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[607-:32] + 6) >= 7 ? hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[607-:32] + 0 : 8 - (hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[607-:32] + 6))];
	assign axi_aw_o[aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_AddrWidth + (29 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 5))-:((aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_AddrWidth + (29 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 5))) >= (35 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 0)) ? ((aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_AddrWidth + (29 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 5))) - (35 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 0))) + 1 : ((35 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 0)) - (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_AddrWidth + (29 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 5)))) + 1)] = req_i[hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[639-:32] + (11 + (hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[607-:32] + 6))-:((hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[639-:32] + (11 + (hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[607-:32] + 6))) >= (11 + (hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[607-:32] + 7)) ? ((hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[639-:32] + (11 + (hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[607-:32] + 6))) - (11 + (hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[607-:32] + 7))) + 1 : ((11 + (hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[607-:32] + 7)) - (hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[639-:32] + (11 + (hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[607-:32] + 6)))) + 1)];
	assign axi_aw_o[29 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 5)-:((29 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 5)) >= (27 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 0)) ? ((29 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 5)) - (27 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 0))) + 1 : ((27 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 0)) - (29 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 5))) + 1)] = req_i[11 + (hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[607-:32] + 6)-:((11 + (hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[607-:32] + 6)) >= (3 + (hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[607-:32] + 7)) ? ((11 + (hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[607-:32] + 6)) - (3 + (hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[607-:32] + 7))) + 1 : ((3 + (hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[607-:32] + 7)) - (11 + (hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[607-:32] + 6))) + 1)];
	assign axi_aw_o[17 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 9)-:((17 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 9)) >= (24 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 0)) ? ((17 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 9)) - (24 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 0))) + 1 : ((24 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 0)) - (17 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 9))) + 1)] = req_i[3 + (hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[607-:32] + 6)-:((3 + (hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[607-:32] + 6)) >= (hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[607-:32] + 7) ? ((3 + (hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[607-:32] + 6)) - (hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[607-:32] + 7)) + 1 : ((hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[607-:32] + 7) - (3 + (hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[607-:32] + 6))) + 1)];
	localparam axi_pkg_BURST_INCR = 2'b01;
	assign axi_aw_o[18 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 5)-:((18 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 5)) >= (22 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 0)) ? ((18 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 5)) - (22 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 0))) + 1 : ((22 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 0)) - (18 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 5))) + 1)] = axi_pkg_BURST_INCR;
	assign axi_aw_o[12 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 9)] = lock;
	assign axi_aw_o[15 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 5)-:((15 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 5)) >= (17 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 0)) ? ((15 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 5)) - (17 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 0))) + 1 : ((17 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 0)) - (15 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 5))) + 1)] = cache;
	assign axi_aw_o[7 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 9)-:((7 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 9)) >= (14 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 0)) ? ((7 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 9)) - (14 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 0))) + 1 : ((14 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 0)) - (7 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 9))) + 1)] = 1'sb0;
	assign axi_aw_o[8 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 5)-:((8 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 5)) >= (10 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 0)) ? ((8 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 5)) - (10 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 0))) + 1 : ((10 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 0)) - (8 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 5))) + 1)] = 1'sb0;
	assign axi_aw_o[aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 9-:((aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 9) >= (6 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 0)) ? ((aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 9) - (6 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 0))) + 1 : ((6 + (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 0)) - (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 9)) + 1)] = 1'sb0;
	assign axi_aw_o[aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 5-:((aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 5) >= (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 0) ? ((aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 5) - (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 0)) + 1 : ((aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 0) - (aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth + 5)) + 1)] = atop;
	assign axi_aw_o[aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth - 1-:aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_axi_aw_chan_t_ariane_axi_UserWidth] = 1'sb0;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_write.sv:135:5
	assign req_data_ready_o = axi_w_ready_i;
	assign axi_w_valid_o = req_data_valid_i;
	assign axi_w_o[w_chan_t_axi_w_chan_t_axi_w_chan_t_axi_w_chan_t_ariane_axi_DataWidth + (w_chan_t_axi_w_chan_t_axi_w_chan_t_axi_w_chan_t_ariane_axi_StrbWidth + (w_chan_t_axi_w_chan_t_axi_w_chan_t_axi_w_chan_t_ariane_axi_UserWidth + 0))-:((w_chan_t_axi_w_chan_t_axi_w_chan_t_axi_w_chan_t_ariane_axi_DataWidth + (w_chan_t_axi_w_chan_t_axi_w_chan_t_axi_w_chan_t_ariane_axi_StrbWidth + (w_chan_t_axi_w_chan_t_axi_w_chan_t_axi_w_chan_t_ariane_axi_UserWidth + 0))) >= (w_chan_t_axi_w_chan_t_axi_w_chan_t_axi_w_chan_t_ariane_axi_StrbWidth + (1 + (w_chan_t_axi_w_chan_t_axi_w_chan_t_axi_w_chan_t_ariane_axi_UserWidth + 0))) ? ((w_chan_t_axi_w_chan_t_axi_w_chan_t_axi_w_chan_t_ariane_axi_DataWidth + (w_chan_t_axi_w_chan_t_axi_w_chan_t_axi_w_chan_t_ariane_axi_StrbWidth + (w_chan_t_axi_w_chan_t_axi_w_chan_t_axi_w_chan_t_ariane_axi_UserWidth + 0))) - (w_chan_t_axi_w_chan_t_axi_w_chan_t_axi_w_chan_t_ariane_axi_StrbWidth + (1 + (w_chan_t_axi_w_chan_t_axi_w_chan_t_axi_w_chan_t_ariane_axi_UserWidth + 0)))) + 1 : ((w_chan_t_axi_w_chan_t_axi_w_chan_t_axi_w_chan_t_ariane_axi_StrbWidth + (1 + (w_chan_t_axi_w_chan_t_axi_w_chan_t_axi_w_chan_t_ariane_axi_UserWidth + 0))) - (w_chan_t_axi_w_chan_t_axi_w_chan_t_axi_w_chan_t_ariane_axi_DataWidth + (w_chan_t_axi_w_chan_t_axi_w_chan_t_axi_w_chan_t_ariane_axi_StrbWidth + (w_chan_t_axi_w_chan_t_axi_w_chan_t_axi_w_chan_t_ariane_axi_UserWidth + 0)))) + 1)] = req_data_i[hpdcache_mem_req_w_t_hpdcache_mem_req_w_t_HPDcacheCfg[575-:32] + ((hpdcache_mem_req_w_t_hpdcache_mem_req_w_t_HPDcacheCfg[575-:32] / 8) + 0)-:((hpdcache_mem_req_w_t_hpdcache_mem_req_w_t_HPDcacheCfg[575-:32] + ((hpdcache_mem_req_w_t_hpdcache_mem_req_w_t_HPDcacheCfg[575-:32] / 8) + 0)) >= ((hpdcache_mem_req_w_t_hpdcache_mem_req_w_t_HPDcacheCfg[575-:32] / 8) + 1) ? ((hpdcache_mem_req_w_t_hpdcache_mem_req_w_t_HPDcacheCfg[575-:32] + ((hpdcache_mem_req_w_t_hpdcache_mem_req_w_t_HPDcacheCfg[575-:32] / 8) + 0)) - ((hpdcache_mem_req_w_t_hpdcache_mem_req_w_t_HPDcacheCfg[575-:32] / 8) + 1)) + 1 : (((hpdcache_mem_req_w_t_hpdcache_mem_req_w_t_HPDcacheCfg[575-:32] / 8) + 1) - (hpdcache_mem_req_w_t_hpdcache_mem_req_w_t_HPDcacheCfg[575-:32] + ((hpdcache_mem_req_w_t_hpdcache_mem_req_w_t_HPDcacheCfg[575-:32] / 8) + 0))) + 1)];
	assign axi_w_o[w_chan_t_axi_w_chan_t_axi_w_chan_t_axi_w_chan_t_ariane_axi_StrbWidth + (w_chan_t_axi_w_chan_t_axi_w_chan_t_axi_w_chan_t_ariane_axi_UserWidth + 0)-:((w_chan_t_axi_w_chan_t_axi_w_chan_t_axi_w_chan_t_ariane_axi_StrbWidth + (w_chan_t_axi_w_chan_t_axi_w_chan_t_axi_w_chan_t_ariane_axi_UserWidth + 0)) >= (1 + (w_chan_t_axi_w_chan_t_axi_w_chan_t_axi_w_chan_t_ariane_axi_UserWidth + 0)) ? ((w_chan_t_axi_w_chan_t_axi_w_chan_t_axi_w_chan_t_ariane_axi_StrbWidth + (w_chan_t_axi_w_chan_t_axi_w_chan_t_axi_w_chan_t_ariane_axi_UserWidth + 0)) - (1 + (w_chan_t_axi_w_chan_t_axi_w_chan_t_axi_w_chan_t_ariane_axi_UserWidth + 0))) + 1 : ((1 + (w_chan_t_axi_w_chan_t_axi_w_chan_t_axi_w_chan_t_ariane_axi_UserWidth + 0)) - (w_chan_t_axi_w_chan_t_axi_w_chan_t_axi_w_chan_t_ariane_axi_StrbWidth + (w_chan_t_axi_w_chan_t_axi_w_chan_t_axi_w_chan_t_ariane_axi_UserWidth + 0))) + 1)] = req_data_i[(hpdcache_mem_req_w_t_hpdcache_mem_req_w_t_HPDcacheCfg[575-:32] / 8) + 0-:(((hpdcache_mem_req_w_t_hpdcache_mem_req_w_t_HPDcacheCfg[575-:32] / 8) + 0) >= 1 ? (hpdcache_mem_req_w_t_hpdcache_mem_req_w_t_HPDcacheCfg[575-:32] / 8) + 0 : 2 - ((hpdcache_mem_req_w_t_hpdcache_mem_req_w_t_HPDcacheCfg[575-:32] / 8) + 0))];
	assign axi_w_o[w_chan_t_axi_w_chan_t_axi_w_chan_t_axi_w_chan_t_ariane_axi_UserWidth + 0] = req_data_i[0];
	assign axi_w_o[w_chan_t_axi_w_chan_t_axi_w_chan_t_axi_w_chan_t_ariane_axi_UserWidth - 1-:w_chan_t_axi_w_chan_t_axi_w_chan_t_axi_w_chan_t_ariane_axi_UserWidth] = 1'sb0;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_write.sv:142:5
	assign axi_b_ready_o = resp_ready_i;
	assign resp_valid_o = axi_b_valid_i;
	assign resp_o[hpdcache_mem_resp_w_t_hpdcache_mem_resp_w_t_HPDcacheCfg[607-:32] + 1-:((hpdcache_mem_resp_w_t_hpdcache_mem_resp_w_t_HPDcacheCfg[607-:32] + 1) >= (hpdcache_mem_resp_w_t_hpdcache_mem_resp_w_t_HPDcacheCfg[607-:32] + 0) ? ((hpdcache_mem_resp_w_t_hpdcache_mem_resp_w_t_HPDcacheCfg[607-:32] + 1) - (hpdcache_mem_resp_w_t_hpdcache_mem_resp_w_t_HPDcacheCfg[607-:32] + 0)) + 1 : ((hpdcache_mem_resp_w_t_hpdcache_mem_resp_w_t_HPDcacheCfg[607-:32] + 0) - (hpdcache_mem_resp_w_t_hpdcache_mem_resp_w_t_HPDcacheCfg[607-:32] + 1)) + 1)] = resp;
	assign resp_o[hpdcache_mem_resp_w_t_hpdcache_mem_resp_w_t_HPDcacheCfg[607-:32] - 1-:hpdcache_mem_resp_w_t_hpdcache_mem_resp_w_t_HPDcacheCfg[607-:32]] = axi_b_i[b_chan_t_axi_b_chan_t_axi_b_chan_t_CVA6Cfg[9119 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9119 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9119 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9119 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (b_chan_t_axi_b_chan_t_axi_b_chan_t_CVA6Cfg[9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 1)-:((b_chan_t_axi_b_chan_t_axi_b_chan_t_CVA6Cfg[9119 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9119 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9119 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9119 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (b_chan_t_axi_b_chan_t_axi_b_chan_t_CVA6Cfg[9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 1)) >= (2 + (b_chan_t_axi_b_chan_t_axi_b_chan_t_CVA6Cfg[9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0)) ? ((b_chan_t_axi_b_chan_t_axi_b_chan_t_CVA6Cfg[9119 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9119 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9119 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9119 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (b_chan_t_axi_b_chan_t_axi_b_chan_t_CVA6Cfg[9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 1)) - (2 + (b_chan_t_axi_b_chan_t_axi_b_chan_t_CVA6Cfg[9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0))) + 1 : ((2 + (b_chan_t_axi_b_chan_t_axi_b_chan_t_CVA6Cfg[9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0)) - (b_chan_t_axi_b_chan_t_axi_b_chan_t_CVA6Cfg[9119 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9119 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9119 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9119 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (b_chan_t_axi_b_chan_t_axi_b_chan_t_CVA6Cfg[9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 1))) + 1)];
	localparam axi_pkg_RESP_EXOKAY = 2'b01;
	assign resp_o[hpdcache_mem_resp_w_t_hpdcache_mem_resp_w_t_HPDcacheCfg[607-:32] + 2] = axi_b_i[b_chan_t_axi_b_chan_t_axi_b_chan_t_CVA6Cfg[9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 1-:((b_chan_t_axi_b_chan_t_axi_b_chan_t_CVA6Cfg[9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 1) >= (b_chan_t_axi_b_chan_t_axi_b_chan_t_CVA6Cfg[9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0) ? ((b_chan_t_axi_b_chan_t_axi_b_chan_t_CVA6Cfg[9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 1) - (b_chan_t_axi_b_chan_t_axi_b_chan_t_CVA6Cfg[9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0)) + 1 : ((b_chan_t_axi_b_chan_t_axi_b_chan_t_CVA6Cfg[9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0) - (b_chan_t_axi_b_chan_t_axi_b_chan_t_CVA6Cfg[9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9055 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9087 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + ((b_chan_t_axi_b_chan_t_axi_b_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 1)) + 1)] == axi_pkg_RESP_EXOKAY;
	initial _sv2v_0 = 0;
endmodule
