module hpdcache_ctrl_9FAF1_89982 (
	clk_i,
	rst_ni,
	core_req_valid_i,
	core_req_ready_o,
	core_req_i,
	core_req_abort_i,
	core_req_tag_i,
	core_req_pma_i,
	core_rsp_valid_o,
	core_rsp_o,
	wbuf_flush_i,
	cachedir_hit_o,
	miss_mshr_check_o,
	miss_mshr_check_offset_o,
	miss_mshr_check_nline_o,
	miss_mshr_alloc_o,
	miss_mshr_alloc_cs_o,
	miss_mshr_alloc_ready_i,
	miss_mshr_alloc_full_i,
	miss_mshr_alloc_nline_o,
	miss_mshr_alloc_tid_o,
	miss_mshr_alloc_sid_o,
	miss_mshr_alloc_word_o,
	miss_mshr_alloc_need_rsp_o,
	miss_mshr_alloc_is_prefetch_o,
	miss_mshr_hit_i,
	refill_req_valid_i,
	refill_req_ready_o,
	refill_busy_i,
	refill_sel_victim_i,
	refill_updt_plru_i,
	refill_set_i,
	refill_dir_entry_i,
	refill_victim_way_o,
	refill_victim_way_i,
	refill_write_dir_i,
	refill_write_data_i,
	refill_word_i,
	refill_data_i,
	refill_core_rsp_valid_i,
	refill_core_rsp_i,
	refill_nline_i,
	refill_updt_rtab_i,
	inval_check_dir_i,
	inval_write_dir_i,
	inval_nline_i,
	inval_hit_o,
	wbuf_empty_i,
	wbuf_flush_all_o,
	wbuf_write_o,
	wbuf_write_ready_i,
	wbuf_write_addr_o,
	wbuf_write_data_o,
	wbuf_write_be_o,
	wbuf_write_uncacheable_o,
	wbuf_read_hit_i,
	wbuf_read_flush_hit_o,
	wbuf_rtab_addr_o,
	wbuf_rtab_is_read_o,
	wbuf_rtab_hit_open_i,
	wbuf_rtab_hit_pend_i,
	wbuf_rtab_hit_sent_i,
	wbuf_rtab_not_ready_i,
	uc_busy_i,
	uc_lrsc_snoop_o,
	uc_lrsc_snoop_addr_o,
	uc_lrsc_snoop_size_o,
	uc_req_valid_o,
	uc_req_op_o,
	uc_req_addr_o,
	uc_req_size_o,
	uc_req_data_o,
	uc_req_be_o,
	uc_req_uc_o,
	uc_req_sid_o,
	uc_req_tid_o,
	uc_req_need_rsp_o,
	uc_wbuf_flush_all_i,
	uc_dir_amo_match_i,
	uc_dir_amo_match_set_i,
	uc_dir_amo_match_tag_i,
	uc_dir_amo_update_plru_i,
	uc_dir_amo_hit_way_o,
	uc_data_amo_write_i,
	uc_data_amo_write_enable_i,
	uc_data_amo_write_set_i,
	uc_data_amo_write_size_i,
	uc_data_amo_write_word_i,
	uc_data_amo_write_data_i,
	uc_data_amo_write_be_i,
	uc_core_rsp_ready_o,
	uc_core_rsp_valid_i,
	uc_core_rsp_i,
	cmo_busy_i,
	cmo_wait_i,
	cmo_req_valid_o,
	cmo_req_op_o,
	cmo_req_addr_o,
	cmo_req_wdata_o,
	cmo_wbuf_flush_all_i,
	cmo_dir_check_i,
	cmo_dir_check_set_i,
	cmo_dir_check_tag_i,
	cmo_dir_check_hit_way_o,
	cmo_dir_inval_i,
	cmo_dir_inval_set_i,
	cmo_dir_inval_way_i,
	rtab_empty_o,
	ctrl_empty_o,
	cfg_enable_i,
	cfg_rtab_single_entry_i,
	evt_cache_write_miss_o,
	evt_cache_read_miss_o,
	evt_uncached_req_o,
	evt_cmo_req_o,
	evt_write_req_o,
	evt_read_req_o,
	evt_prefetch_req_o,
	evt_req_on_hold_o,
	evt_rtab_rollback_o,
	evt_stall_refill_o,
	evt_stall_o
);
	// removed localparam type hpdcache_data_be_t_hpdcache_data_be_t_hpdcache_data_be_t_HPDcacheCfg_type
	parameter [1349:0] hpdcache_data_be_t_hpdcache_data_be_t_hpdcache_data_be_t_HPDcacheCfg = 0;
	// removed localparam type hpdcache_data_word_t_hpdcache_data_word_t_hpdcache_data_word_t_HPDcacheCfg_type
	parameter [1349:0] hpdcache_data_word_t_hpdcache_data_word_t_hpdcache_data_word_t_HPDcacheCfg = 0;
	// removed localparam type hpdcache_dir_entry_t_hpdcache_tag_t_hpdcache_tag_t_HPDcacheCfg_type
	parameter [1349:0] hpdcache_dir_entry_t_hpdcache_tag_t_hpdcache_tag_t_HPDcacheCfg = 0;
	// removed localparam type hpdcache_nline_t_HPDcacheCfg_type
	parameter [1349:0] hpdcache_nline_t_HPDcacheCfg = 0;
	// removed localparam type hpdcache_refill_be_t_HPDcacheCfg_type
	// removed localparam type hpdcache_refill_be_t_hpdcache_data_be_t_hpdcache_data_be_t_HPDcacheCfg_type
	parameter [1349:0] hpdcache_refill_be_t_HPDcacheCfg = 0;
	parameter [1349:0] hpdcache_refill_be_t_hpdcache_data_be_t_hpdcache_data_be_t_HPDcacheCfg = 0;
	// removed localparam type hpdcache_refill_data_t_HPDcacheCfg_type
	// removed localparam type hpdcache_refill_data_t_hpdcache_data_word_t_hpdcache_data_word_t_HPDcacheCfg_type
	parameter [1349:0] hpdcache_refill_data_t_HPDcacheCfg = 0;
	parameter [1349:0] hpdcache_refill_data_t_hpdcache_data_word_t_hpdcache_data_word_t_HPDcacheCfg = 0;
	// removed localparam type hpdcache_req_addr_t_HPDcacheCfg_type
	parameter [1349:0] hpdcache_req_addr_t_HPDcacheCfg = 0;
	// removed localparam type hpdcache_req_be_t_hpdcache_req_be_t_hpdcache_req_be_t_HPDcacheCfg_type
	parameter [1349:0] hpdcache_req_be_t_hpdcache_req_be_t_hpdcache_req_be_t_HPDcacheCfg = 0;
	// removed localparam type hpdcache_req_data_t_hpdcache_req_data_t_hpdcache_req_data_t_HPDcacheCfg_type
	parameter [1349:0] hpdcache_req_data_t_hpdcache_req_data_t_hpdcache_req_data_t_HPDcacheCfg = 0;
	// removed localparam type hpdcache_req_offset_t_hpdcache_req_offset_t_hpdcache_req_offset_t_HPDcacheCfg_type
	parameter [1349:0] hpdcache_req_offset_t_hpdcache_req_offset_t_hpdcache_req_offset_t_HPDcacheCfg = 0;
	// removed localparam type hpdcache_req_sid_t_hpdcache_req_sid_t_hpdcache_req_sid_t_HPDcacheCfg_type
	parameter [1349:0] hpdcache_req_sid_t_hpdcache_req_sid_t_hpdcache_req_sid_t_HPDcacheCfg = 0;
	// removed localparam type hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg_type
	parameter [1349:0] hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg = 0;
	// removed localparam type hpdcache_req_tid_t_hpdcache_req_tid_t_hpdcache_req_tid_t_HPDcacheCfg_type
	parameter [1349:0] hpdcache_req_tid_t_hpdcache_req_tid_t_hpdcache_req_tid_t_HPDcacheCfg = 0;
	// removed localparam type hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg_type
	parameter [1349:0] hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg = 0;
	// removed localparam type hpdcache_set_t_HPDcacheCfg_type
	parameter [1349:0] hpdcache_set_t_HPDcacheCfg = 0;
	// removed localparam type hpdcache_tag_t_hpdcache_tag_t_hpdcache_tag_t_HPDcacheCfg_type
	parameter [1349:0] hpdcache_tag_t_hpdcache_tag_t_hpdcache_tag_t_HPDcacheCfg = 0;
	// removed localparam type hpdcache_way_vector_t_HPDcacheCfg_type
	parameter [1349:0] hpdcache_way_vector_t_HPDcacheCfg = 0;
	// removed localparam type hpdcache_word_t_HPDcacheCfg_type
	parameter [1349:0] hpdcache_word_t_HPDcacheCfg = 0;
	// removed localparam type wbuf_addr_t_HPDcacheCfg_type
	parameter [1349:0] wbuf_addr_t_HPDcacheCfg = 0;
	// removed localparam type wbuf_be_t_hpdcache_req_be_t_hpdcache_req_be_t_HPDcacheCfg_type
	parameter [1349:0] wbuf_be_t_hpdcache_req_be_t_hpdcache_req_be_t_HPDcacheCfg = 0;
	// removed localparam type wbuf_data_t_hpdcache_req_data_t_hpdcache_req_data_t_HPDcacheCfg_type
	parameter [1349:0] wbuf_data_t_hpdcache_req_data_t_hpdcache_req_data_t_HPDcacheCfg = 0;
	// removed import hpdcache_pkg::*;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:35:15
	// removed localparam type hpdcache_pkg_hpdcache_victim_sel_policy_t
	// removed localparam type hpdcache_pkg_hpdcache_user_cfg_t
	// removed localparam type hpdcache_pkg_hpdcache_cfg_t
	parameter [1349:0] HPDcacheCfg = 1'sb0;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:37:20
	// removed localparam type hpdcache_nline_t
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:38:20
	// removed localparam type hpdcache_tag_t
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:39:20
	// removed localparam type hpdcache_set_t
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:40:20
	// removed localparam type hpdcache_word_t
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:41:20
	// removed localparam type hpdcache_data_word_t
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:42:20
	// removed localparam type hpdcache_data_be_t
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:43:20
	// removed localparam type hpdcache_dir_entry_t
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:44:20
	// removed localparam type hpdcache_way_vector_t
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:46:20
	// removed localparam type wbuf_addr_t
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:47:20
	// removed localparam type wbuf_data_t
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:48:20
	// removed localparam type wbuf_be_t
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:50:20
	// removed localparam type hpdcache_refill_data_t
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:51:20
	// removed localparam type hpdcache_refill_be_t
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:53:20
	// removed localparam type hpdcache_req_addr_t
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:54:20
	// removed localparam type hpdcache_req_offset_t
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:55:20
	// removed localparam type hpdcache_req_tid_t
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:56:20
	// removed localparam type hpdcache_req_sid_t
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:57:20
	// removed localparam type hpdcache_req_data_t
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:58:20
	// removed localparam type hpdcache_req_be_t
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:60:20
	// removed localparam type hpdcache_req_t
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:61:20
	// removed localparam type hpdcache_rsp_t
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:68:5
	input wire clk_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:69:5
	input wire rst_ni;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:72:5
	input wire core_req_valid_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:73:5
	output wire core_req_ready_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:74:5
	input wire [((((((((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1:0] core_req_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:75:5
	input wire core_req_abort_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:76:5
	input wire [hpdcache_tag_t_hpdcache_tag_t_hpdcache_tag_t_HPDcacheCfg[351-:32] - 1:0] core_req_tag_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:77:5
	// removed localparam type hpdcache_pkg_hpdcache_pma_t
	input wire [1:0] core_req_pma_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:80:5
	output wire core_rsp_valid_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:81:5
	output wire [(((hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1157-:32] * hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1285-:32]) + hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32]) + hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32]) + 1:0] core_rsp_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:84:5
	input wire wbuf_flush_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:87:5
	output wire cachedir_hit_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:90:5
	output wire miss_mshr_check_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:91:5
	output wire [hpdcache_req_offset_t_hpdcache_req_offset_t_hpdcache_req_offset_t_HPDcacheCfg[287-:32] - 1:0] miss_mshr_check_offset_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:92:5
	output wire [hpdcache_nline_t_HPDcacheCfg[383-:32] - 1:0] miss_mshr_check_nline_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:93:5
	output wire miss_mshr_alloc_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:94:5
	output wire miss_mshr_alloc_cs_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:95:5
	input wire miss_mshr_alloc_ready_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:96:5
	input wire miss_mshr_alloc_full_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:97:5
	output wire [hpdcache_nline_t_HPDcacheCfg[383-:32] - 1:0] miss_mshr_alloc_nline_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:98:5
	output wire [hpdcache_req_tid_t_hpdcache_req_tid_t_hpdcache_req_tid_t_HPDcacheCfg[1125-:32] - 1:0] miss_mshr_alloc_tid_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:99:5
	output wire [hpdcache_req_sid_t_hpdcache_req_sid_t_hpdcache_req_sid_t_HPDcacheCfg[1093-:32] - 1:0] miss_mshr_alloc_sid_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:100:5
	output wire [hpdcache_word_t_HPDcacheCfg[511-:32] - 1:0] miss_mshr_alloc_word_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:101:5
	output wire miss_mshr_alloc_need_rsp_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:102:5
	output wire miss_mshr_alloc_is_prefetch_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:103:5
	input wire miss_mshr_hit_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:106:5
	input wire refill_req_valid_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:107:5
	output wire refill_req_ready_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:108:5
	input wire refill_busy_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:109:5
	input wire refill_sel_victim_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:110:5
	input wire refill_updt_plru_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:111:5
	input wire [hpdcache_set_t_HPDcacheCfg[415-:32] - 1:0] refill_set_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:112:5
	input wire [(1 + hpdcache_dir_entry_t_hpdcache_tag_t_hpdcache_tag_t_HPDcacheCfg[351-:32]) + 0:0] refill_dir_entry_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:113:5
	output wire [hpdcache_way_vector_t_HPDcacheCfg[1221-:32] - 1:0] refill_victim_way_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:114:5
	input wire [hpdcache_way_vector_t_HPDcacheCfg[1221-:32] - 1:0] refill_victim_way_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:115:5
	input wire refill_write_dir_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:116:5
	input wire refill_write_data_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:117:5
	input wire [hpdcache_word_t_HPDcacheCfg[511-:32] - 1:0] refill_word_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:118:5
	input wire [(hpdcache_refill_data_t_HPDcacheCfg[995-:32] * hpdcache_refill_data_t_hpdcache_data_word_t_hpdcache_data_word_t_HPDcacheCfg[1285-:32]) - 1:0] refill_data_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:119:5
	input wire refill_core_rsp_valid_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:120:5
	input wire [(((hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1157-:32] * hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1285-:32]) + hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32]) + hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32]) + 1:0] refill_core_rsp_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:121:5
	input wire [hpdcache_nline_t_HPDcacheCfg[383-:32] - 1:0] refill_nline_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:122:5
	input wire refill_updt_rtab_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:125:5
	input wire inval_check_dir_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:126:5
	input wire inval_write_dir_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:127:5
	input wire [hpdcache_nline_t_HPDcacheCfg[383-:32] - 1:0] inval_nline_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:128:5
	output wire inval_hit_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:131:5
	input wire wbuf_empty_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:132:5
	output wire wbuf_flush_all_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:133:5
	output wire wbuf_write_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:134:5
	input wire wbuf_write_ready_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:135:5
	output wire [wbuf_addr_t_HPDcacheCfg[1317-:32] - 1:0] wbuf_write_addr_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:136:5
	output wire [(wbuf_data_t_hpdcache_req_data_t_hpdcache_req_data_t_HPDcacheCfg[1157-:32] * wbuf_data_t_hpdcache_req_data_t_hpdcache_req_data_t_HPDcacheCfg[1285-:32]) - 1:0] wbuf_write_data_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:137:5
	output wire [(wbuf_be_t_hpdcache_req_be_t_hpdcache_req_be_t_HPDcacheCfg[1157-:32] * (wbuf_be_t_hpdcache_req_be_t_hpdcache_req_be_t_HPDcacheCfg[1285-:32] / 8)) - 1:0] wbuf_write_be_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:138:5
	output wire wbuf_write_uncacheable_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:139:5
	input wire wbuf_read_hit_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:140:5
	output wire wbuf_read_flush_hit_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:141:5
	output wire [hpdcache_req_addr_t_HPDcacheCfg[1317-:32] - 1:0] wbuf_rtab_addr_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:142:5
	output wire wbuf_rtab_is_read_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:143:5
	input wire wbuf_rtab_hit_open_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:144:5
	input wire wbuf_rtab_hit_pend_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:145:5
	input wire wbuf_rtab_hit_sent_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:146:5
	input wire wbuf_rtab_not_ready_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:149:5
	input wire uc_busy_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:150:5
	output wire uc_lrsc_snoop_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:151:5
	output wire [hpdcache_req_addr_t_HPDcacheCfg[1317-:32] - 1:0] uc_lrsc_snoop_addr_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:152:5
	// removed localparam type hpdcache_pkg_hpdcache_req_size_t
	output wire [2:0] uc_lrsc_snoop_size_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:153:5
	output wire uc_req_valid_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:154:5
	// removed localparam type hpdcache_pkg_hpdcache_uc_op_t
	output wire [12:0] uc_req_op_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:155:5
	output wire [hpdcache_req_addr_t_HPDcacheCfg[1317-:32] - 1:0] uc_req_addr_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:156:5
	output wire [2:0] uc_req_size_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:157:5
	output wire [(hpdcache_req_data_t_hpdcache_req_data_t_hpdcache_req_data_t_HPDcacheCfg[1157-:32] * hpdcache_req_data_t_hpdcache_req_data_t_hpdcache_req_data_t_HPDcacheCfg[1285-:32]) - 1:0] uc_req_data_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:158:5
	output wire [(hpdcache_req_be_t_hpdcache_req_be_t_hpdcache_req_be_t_HPDcacheCfg[1157-:32] * (hpdcache_req_be_t_hpdcache_req_be_t_hpdcache_req_be_t_HPDcacheCfg[1285-:32] / 8)) - 1:0] uc_req_be_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:159:5
	output wire uc_req_uc_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:160:5
	output wire [hpdcache_req_sid_t_hpdcache_req_sid_t_hpdcache_req_sid_t_HPDcacheCfg[1093-:32] - 1:0] uc_req_sid_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:161:5
	output wire [hpdcache_req_tid_t_hpdcache_req_tid_t_hpdcache_req_tid_t_HPDcacheCfg[1125-:32] - 1:0] uc_req_tid_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:162:5
	output wire uc_req_need_rsp_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:163:5
	input wire uc_wbuf_flush_all_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:164:5
	input wire uc_dir_amo_match_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:165:5
	input wire [hpdcache_set_t_HPDcacheCfg[415-:32] - 1:0] uc_dir_amo_match_set_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:166:5
	input wire [hpdcache_tag_t_hpdcache_tag_t_hpdcache_tag_t_HPDcacheCfg[351-:32] - 1:0] uc_dir_amo_match_tag_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:167:5
	input wire uc_dir_amo_update_plru_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:168:5
	output wire [hpdcache_way_vector_t_HPDcacheCfg[1221-:32] - 1:0] uc_dir_amo_hit_way_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:169:5
	input wire uc_data_amo_write_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:170:5
	input wire uc_data_amo_write_enable_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:171:5
	input wire [hpdcache_set_t_HPDcacheCfg[415-:32] - 1:0] uc_data_amo_write_set_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:172:5
	input wire [2:0] uc_data_amo_write_size_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:173:5
	input wire [hpdcache_word_t_HPDcacheCfg[511-:32] - 1:0] uc_data_amo_write_word_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:174:5
	input wire [(hpdcache_req_data_t_hpdcache_req_data_t_hpdcache_req_data_t_HPDcacheCfg[1157-:32] * hpdcache_req_data_t_hpdcache_req_data_t_hpdcache_req_data_t_HPDcacheCfg[1285-:32]) - 1:0] uc_data_amo_write_data_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:175:5
	input wire [(hpdcache_req_be_t_hpdcache_req_be_t_hpdcache_req_be_t_HPDcacheCfg[1157-:32] * (hpdcache_req_be_t_hpdcache_req_be_t_hpdcache_req_be_t_HPDcacheCfg[1285-:32] / 8)) - 1:0] uc_data_amo_write_be_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:176:5
	output wire uc_core_rsp_ready_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:177:5
	input wire uc_core_rsp_valid_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:178:5
	input wire [(((hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1157-:32] * hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1285-:32]) + hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32]) + hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32]) + 1:0] uc_core_rsp_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:181:5
	input wire cmo_busy_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:182:5
	input wire cmo_wait_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:183:5
	output wire cmo_req_valid_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:184:5
	// removed localparam type hpdcache_pkg_hpdcache_cmoh_op_t
	output wire [3:0] cmo_req_op_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:185:5
	output wire [hpdcache_req_addr_t_HPDcacheCfg[1317-:32] - 1:0] cmo_req_addr_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:186:5
	output wire [(hpdcache_req_data_t_hpdcache_req_data_t_hpdcache_req_data_t_HPDcacheCfg[1157-:32] * hpdcache_req_data_t_hpdcache_req_data_t_hpdcache_req_data_t_HPDcacheCfg[1285-:32]) - 1:0] cmo_req_wdata_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:187:5
	input wire cmo_wbuf_flush_all_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:188:5
	input wire cmo_dir_check_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:189:5
	input wire [hpdcache_set_t_HPDcacheCfg[415-:32] - 1:0] cmo_dir_check_set_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:190:5
	input wire [hpdcache_tag_t_hpdcache_tag_t_hpdcache_tag_t_HPDcacheCfg[351-:32] - 1:0] cmo_dir_check_tag_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:191:5
	output wire [hpdcache_way_vector_t_HPDcacheCfg[1221-:32] - 1:0] cmo_dir_check_hit_way_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:192:5
	input wire cmo_dir_inval_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:193:5
	input wire [hpdcache_set_t_HPDcacheCfg[415-:32] - 1:0] cmo_dir_inval_set_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:194:5
	input wire [hpdcache_way_vector_t_HPDcacheCfg[1221-:32] - 1:0] cmo_dir_inval_way_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:196:5
	output wire rtab_empty_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:197:5
	output wire ctrl_empty_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:200:5
	input wire cfg_enable_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:201:5
	input wire cfg_rtab_single_entry_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:204:5
	output wire evt_cache_write_miss_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:205:5
	output wire evt_cache_read_miss_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:206:5
	output wire evt_uncached_req_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:207:5
	output wire evt_cmo_req_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:208:5
	output wire evt_write_req_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:209:5
	output wire evt_read_req_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:210:5
	output wire evt_prefetch_req_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:211:5
	output wire evt_req_on_hold_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:212:5
	output wire evt_rtab_rollback_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:213:5
	output wire evt_stall_refill_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:214:5
	output wire evt_stall_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:220:5
	// removed localparam type rtab_ptr_t
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:225:5
	reg st1_req_valid_q;
	wire st1_req_valid_d;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:226:5
	reg [((((((((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1:0] st1_req_q;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:227:5
	reg st1_req_rtab_q;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:228:5
	reg [$clog2($signed(HPDcacheCfg[671-:32])) - 1:0] st1_rtab_pop_try_ptr_q;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:230:5
	reg st2_req_valid_q;
	wire st2_req_valid_d;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:231:5
	reg st2_req_is_prefetch_q;
	wire st2_req_is_prefetch_d;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:232:5
	reg st2_req_need_rsp_q;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:233:5
	reg [hpdcache_req_addr_t_HPDcacheCfg[1317-:32] - 1:0] st2_req_addr_q;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:234:5
	reg [hpdcache_req_sid_t_hpdcache_req_sid_t_hpdcache_req_sid_t_HPDcacheCfg[1093-:32] - 1:0] st2_req_sid_q;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:235:5
	reg [hpdcache_req_tid_t_hpdcache_req_tid_t_hpdcache_req_tid_t_HPDcacheCfg[1125-:32] - 1:0] st2_req_tid_q;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:240:5
	wire [((((((((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1:0] st0_req;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:241:5
	wire st0_req_is_uncacheable;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:242:5
	wire st0_req_is_load;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:243:5
	wire st0_req_is_store;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:244:5
	wire st0_req_is_amo;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:245:5
	wire st0_req_is_cmo_fence;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:246:5
	wire st0_req_is_cmo_inval;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:247:5
	wire st0_req_is_cmo_prefetch;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:248:5
	wire st0_req_cachedir_read;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:249:5
	wire st0_req_cachedata_read;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:250:5
	wire [hpdcache_set_t_HPDcacheCfg[415-:32] - 1:0] st0_req_set;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:251:5
	wire [hpdcache_word_t_HPDcacheCfg[511-:32] - 1:0] st0_req_word;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:252:5
	wire st0_rtab_pop_try_valid;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:253:5
	wire st0_rtab_pop_try_ready;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:254:5
	wire [((((((((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1:0] st0_rtab_pop_try_req;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:255:5
	wire [$clog2($signed(HPDcacheCfg[671-:32])) - 1:0] st0_rtab_pop_try_ptr;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:257:5
	wire st1_rsp_valid;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:258:5
	wire st1_rsp_aborted;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:259:5
	wire [((((((((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1:0] st1_req;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:260:5
	wire st1_req_abort;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:261:5
	wire st1_req_cachedata_write;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:262:5
	wire st1_req_cachedata_write_enable;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:263:5
	wire [1:0] st1_req_pma;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:264:5
	wire [hpdcache_tag_t_hpdcache_tag_t_hpdcache_tag_t_HPDcacheCfg[351-:32] - 1:0] st1_req_tag;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:265:5
	wire [hpdcache_set_t_HPDcacheCfg[415-:32] - 1:0] st1_req_set;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:266:5
	wire [hpdcache_word_t_HPDcacheCfg[511-:32] - 1:0] st1_req_word;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:267:5
	wire [hpdcache_nline_t_HPDcacheCfg[383-:32] - 1:0] st1_req_nline;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:268:5
	wire [hpdcache_req_addr_t_HPDcacheCfg[1317-:32] - 1:0] st1_req_addr;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:269:5
	wire st1_req_updt_lru;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:270:5
	wire st1_req_is_uncacheable;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:271:5
	wire st1_req_is_load;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:272:5
	wire st1_req_is_store;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:273:5
	wire st1_req_is_amo;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:274:5
	wire st1_req_is_amo_lr;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:275:5
	wire st1_req_is_amo_sc;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:276:5
	wire st1_req_is_amo_swap;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:277:5
	wire st1_req_is_amo_add;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:278:5
	wire st1_req_is_amo_and;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:279:5
	wire st1_req_is_amo_or;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:280:5
	wire st1_req_is_amo_xor;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:281:5
	wire st1_req_is_amo_max;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:282:5
	wire st1_req_is_amo_maxu;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:283:5
	wire st1_req_is_amo_min;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:284:5
	wire st1_req_is_amo_minu;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:285:5
	wire st1_req_is_cmo_inval;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:286:5
	wire st1_req_is_cmo_fence;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:287:5
	wire st1_req_is_cmo_prefetch;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:288:5
	wire [hpdcache_way_vector_t_HPDcacheCfg[1221-:32] - 1:0] st1_dir_hit;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:289:5
	wire [(hpdcache_req_data_t_hpdcache_req_data_t_hpdcache_req_data_t_HPDcacheCfg[1157-:32] * hpdcache_req_data_t_hpdcache_req_data_t_hpdcache_req_data_t_HPDcacheCfg[1285-:32]) - 1:0] st1_read_data;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:290:5
	wire st1_rtab_alloc;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:291:5
	wire st1_rtab_alloc_and_link;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:292:5
	wire st1_rtab_pop_try_commit;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:293:5
	wire st1_rtab_pop_try_rback;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:294:5
	wire st1_rtab_mshr_hit;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:295:5
	wire st1_rtab_mshr_full;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:296:5
	wire st1_rtab_mshr_ready;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:297:5
	wire st1_rtab_wbuf_hit;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:298:5
	wire st1_rtab_wbuf_not_ready;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:299:5
	wire st1_rtab_check;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:300:5
	wire st1_rtab_check_hit;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:302:5
	wire st2_req_we;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:303:5
	wire [hpdcache_word_t_HPDcacheCfg[511-:32] - 1:0] st2_req_word;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:305:5
	wire rtab_full;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:307:5
	wire hpdcache_init_ready;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:313:5
	assign st0_req[hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))-:((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))) >= ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))))) ? ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))))) + 1 : (((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))))) - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))))) + 1)] = (st0_rtab_pop_try_valid ? st0_rtab_pop_try_req[hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))-:((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))) >= ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))))) ? ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))))) + 1 : (((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))))) - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))))) + 1)] : core_req_i[hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))-:((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))) >= ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))))) ? ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))))) + 1 : (((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))))) - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))))) + 1)]);
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:315:5
	assign st0_req[hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1-:((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1) >= 2 ? hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 0 : 3 - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))] = (st0_rtab_pop_try_valid ? st0_rtab_pop_try_req[hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1-:((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1) >= 2 ? hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 0 : 3 - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))] : core_req_i[hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1-:((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1) >= 2 ? hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 0 : 3 - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))]);
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:317:5
	assign st0_req[(hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))-:(((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) >= (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) ? (((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) - (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))))) + 1 : ((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))) + 1)] = (st0_rtab_pop_try_valid ? st0_rtab_pop_try_req[(hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))-:(((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) >= (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) ? (((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) - (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))))) + 1 : ((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))) + 1)] : core_req_i[(hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))-:(((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) >= (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) ? (((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) - (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))))) + 1 : ((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))) + 1)]);
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:319:5
	assign st0_req[4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))-:((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) >= ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) ? ((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) + 1 : (((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) - (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) + 1)] = (st0_rtab_pop_try_valid ? st0_rtab_pop_try_req[4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))-:((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) >= ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) ? ((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) + 1 : (((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) - (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) + 1)] : core_req_i[4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))-:((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) >= ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) ? ((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) + 1 : (((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) - (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) + 1)]);
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:321:5
	assign st0_req[(hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))-:(((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) >= (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))) ? (((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) - (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) + 1 : ((3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) + 1)] = (st0_rtab_pop_try_valid ? st0_rtab_pop_try_req[(hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))-:(((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) >= (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))) ? (((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) - (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) + 1 : ((3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) + 1)] : core_req_i[(hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))-:(((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) >= (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))) ? (((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) - (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) + 1 : ((3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) + 1)]);
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:323:5
	assign st0_req[3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))-:((3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) >= (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) ? ((3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))) + 1 : ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) - (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) + 1)] = (st0_rtab_pop_try_valid ? st0_rtab_pop_try_req[3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))-:((3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) >= (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) ? ((3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))) + 1 : ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) - (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) + 1)] : core_req_i[3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))-:((3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) >= (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) ? ((3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))) + 1 : ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) - (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) + 1)]);
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:325:5
	assign st0_req[hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))-:((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))) >= (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))) ? ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))) - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) + 1 : ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))) - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) + 1)] = (st0_rtab_pop_try_valid ? st0_rtab_pop_try_req[hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))-:((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))) >= (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))) ? ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))) - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) + 1 : ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))) - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) + 1)] : core_req_i[hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))-:((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))) >= (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))) ? ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))) - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) + 1 : ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))) - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) + 1)]);
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:327:5
	assign st0_req[hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))-:((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))) >= (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)) ? ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))) - (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))) + 1 : ((2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)) - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))) + 1)] = (st0_rtab_pop_try_valid ? st0_rtab_pop_try_req[hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))-:((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))) >= (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)) ? ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))) - (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))) + 1 : ((2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)) - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))) + 1)] : core_req_i[hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))-:((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))) >= (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)) ? ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))) - (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))) + 1 : ((2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)) - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))) + 1)]);
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:329:5
	assign st0_req[2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)] = (st0_rtab_pop_try_valid ? st0_rtab_pop_try_req[2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)] : core_req_i[2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)]);
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:331:5
	assign st0_req[1 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)] = (st0_rtab_pop_try_valid ? 1'b1 : core_req_i[1 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)]);
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:333:5
	assign st0_req[1-:2] = (st0_rtab_pop_try_valid ? st0_rtab_pop_try_req[1-:2] : core_req_i[1-:2]);
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:337:5
	assign st0_req_is_uncacheable = ~cfg_enable_i | (st0_req[1 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)] & st0_req[1]);
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:339:5
	// removed localparam type hpdcache_pkg_hpdcache_req_op_t
	function automatic hpdcache_pkg_is_load;
		// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_pkg.sv:97:38
		input reg [3:0] op;
		// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_pkg.sv:98:9
		case (op)
			4'h0: hpdcache_pkg_is_load = 1'b1;
			default: hpdcache_pkg_is_load = 1'b0;
		endcase
	endfunction
	assign st0_req_is_load = hpdcache_pkg_is_load(st0_req[4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))-:((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) >= ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) ? ((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) + 1 : (((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) - (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) + 1)]);
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:340:5
	function automatic hpdcache_pkg_is_store;
		// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_pkg.sv:104:39
		input reg [3:0] op;
		// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_pkg.sv:105:9
		case (op)
			4'h1: hpdcache_pkg_is_store = 1'b1;
			default: hpdcache_pkg_is_store = 1'b0;
		endcase
	endfunction
	assign st0_req_is_store = hpdcache_pkg_is_store(st0_req[4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))-:((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) >= ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) ? ((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) + 1 : (((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) - (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) + 1)]);
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:341:5
	function automatic hpdcache_pkg_is_amo;
		// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_pkg.sv:111:37
		input reg [3:0] op;
		// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_pkg.sv:112:9
		case (op)
			4'h4, 4'h5, 4'h6, 4'h7, 4'h8, 4'h9, 4'ha, 4'hb, 4'hc, 4'hd, 4'he: hpdcache_pkg_is_amo = 1'b1;
			default: hpdcache_pkg_is_amo = 1'b0;
		endcase
	endfunction
	assign st0_req_is_amo = hpdcache_pkg_is_amo(st0_req[4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))-:((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) >= ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) ? ((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) + 1 : (((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) - (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) + 1)]);
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:342:5
	// removed localparam type _sv2v_keep_enum_for_params
	function automatic hpdcache_pkg_is_cmo_fence;
		// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_pkg.sv:241:13
		input reg [3:0] op;
		// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_pkg.sv:242:13
		input reg [2:0] sz;
		// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_pkg.sv:243:9
		case (op)
			4'hf:
				// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_pkg.sv:245:17
				hpdcache_pkg_is_cmo_fence = sz == 3'h0;
			default:
				// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_pkg.sv:248:17
				hpdcache_pkg_is_cmo_fence = 1'b0;
		endcase
	endfunction
	assign st0_req_is_cmo_fence = hpdcache_pkg_is_cmo_fence(st0_req[4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))-:((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) >= ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) ? ((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) + 1 : (((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) - (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) + 1)], st0_req[3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))-:((3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) >= (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) ? ((3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))) + 1 : ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) - (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) + 1)]);
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:343:5
	function automatic hpdcache_pkg_is_cmo_inval;
		// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_pkg.sv:208:13
		input reg [3:0] op;
		// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_pkg.sv:209:13
		input reg [2:0] sz;
		// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_pkg.sv:210:9
		case (op)
			4'hf:
				case (sz)
					3'h2, 3'h3, 3'h4:
						// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_pkg.sv:216:21
						hpdcache_pkg_is_cmo_inval = 1'b1;
					default:
						// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_pkg.sv:219:21
						hpdcache_pkg_is_cmo_inval = 1'b0;
				endcase
			default:
				// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_pkg.sv:223:15
				hpdcache_pkg_is_cmo_inval = 1'b0;
		endcase
	endfunction
	assign st0_req_is_cmo_inval = hpdcache_pkg_is_cmo_inval(st0_req[4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))-:((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) >= ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) ? ((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) + 1 : (((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) - (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) + 1)], st0_req[3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))-:((3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) >= (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) ? ((3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))) + 1 : ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) - (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) + 1)]);
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:344:5
	function automatic hpdcache_pkg_is_cmo_prefetch;
		// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_pkg.sv:254:13
		input reg [3:0] op;
		// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_pkg.sv:255:13
		input reg [2:0] sz;
		// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_pkg.sv:256:9
		case (op)
			4'hf:
				// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_pkg.sv:258:17
				hpdcache_pkg_is_cmo_prefetch = sz == 3'h5;
			default:
				// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_pkg.sv:261:17
				hpdcache_pkg_is_cmo_prefetch = 1'b0;
		endcase
	endfunction
	assign st0_req_is_cmo_prefetch = hpdcache_pkg_is_cmo_prefetch(st0_req[4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))-:((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) >= ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) ? ((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) + 1 : (((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) - (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) + 1)], st0_req[3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))-:((3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) >= (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) ? ((3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))) + 1 : ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) - (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) + 1)]);
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:351:5
	assign st1_req_tag = (st1_req_q[1 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)] ? st1_req_q[hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1-:((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1) >= 2 ? hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 0 : 3 - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))] : core_req_tag_i);
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:352:5
	assign st1_req_pma = (st1_req_q[1 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)] ? st1_req_q[1-:2] : core_req_pma_i);
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:354:5
	assign st1_req[hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))-:((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))) >= ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))))) ? ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))))) + 1 : (((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))))) - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))))) + 1)] = st1_req_q[hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))-:((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))) >= ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))))) ? ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))))) + 1 : (((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))))) - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))))) + 1)];
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:355:5
	assign st1_req[hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1-:((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1) >= 2 ? hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 0 : 3 - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))] = (st1_req_rtab_q ? st1_req_q[hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1-:((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1) >= 2 ? hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 0 : 3 - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))] : st1_req_tag);
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:356:5
	assign st1_req[(hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))-:(((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) >= (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) ? (((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) - (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))))) + 1 : ((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))) + 1)] = st1_req_q[(hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))-:(((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) >= (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) ? (((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) - (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))))) + 1 : ((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))) + 1)];
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:357:5
	assign st1_req[4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))-:((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) >= ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) ? ((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) + 1 : (((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) - (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) + 1)] = st1_req_q[4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))-:((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) >= ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) ? ((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) + 1 : (((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) - (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) + 1)];
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:358:5
	assign st1_req[(hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))-:(((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) >= (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))) ? (((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) - (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) + 1 : ((3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) + 1)] = st1_req_q[(hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))-:(((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) >= (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))) ? (((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) - (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) + 1 : ((3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) + 1)];
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:359:5
	assign st1_req[3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))-:((3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) >= (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) ? ((3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))) + 1 : ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) - (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) + 1)] = st1_req_q[3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))-:((3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) >= (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) ? ((3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))) + 1 : ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) - (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) + 1)];
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:360:5
	assign st1_req[hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))-:((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))) >= (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))) ? ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))) - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) + 1 : ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))) - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) + 1)] = st1_req_q[hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))-:((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))) >= (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))) ? ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))) - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) + 1 : ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))) - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) + 1)];
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:361:5
	assign st1_req[hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))-:((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))) >= (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)) ? ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))) - (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))) + 1 : ((2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)) - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))) + 1)] = st1_req_q[hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))-:((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))) >= (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)) ? ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))) - (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))) + 1 : ((2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)) - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))) + 1)];
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:362:5
	assign st1_req[2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)] = st1_req_q[2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)];
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:363:5
	assign st1_req[1 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)] = st1_req_q[1 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)];
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:364:5
	assign st1_req[1-:2] = (st1_req_rtab_q ? st1_req_q[1-:2] : st1_req_pma);
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:368:5
	assign st1_req_abort = core_req_abort_i & ~st1_req[1 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)];
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:370:5
	assign st1_req_is_uncacheable = ~cfg_enable_i | st1_req[1];
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:371:5
	assign st1_req_is_load = hpdcache_pkg_is_load(st1_req[4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))-:((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) >= ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) ? ((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) + 1 : (((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) - (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) + 1)]);
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:372:5
	assign st1_req_is_store = hpdcache_pkg_is_store(st1_req[4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))-:((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) >= ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) ? ((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) + 1 : (((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) - (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) + 1)]);
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:373:5
	assign st1_req_is_amo = hpdcache_pkg_is_amo(st1_req[4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))-:((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) >= ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) ? ((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) + 1 : (((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) - (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) + 1)]);
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:374:5
	function automatic hpdcache_pkg_is_amo_lr;
		// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_pkg.sv:130:40
		input reg [3:0] op;
		// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_pkg.sv:131:9
		case (op)
			4'h4: hpdcache_pkg_is_amo_lr = 1'b1;
			default: hpdcache_pkg_is_amo_lr = 1'b0;
		endcase
	endfunction
	assign st1_req_is_amo_lr = hpdcache_pkg_is_amo_lr(st1_req[4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))-:((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) >= ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) ? ((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) + 1 : (((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) - (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) + 1)]);
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:375:5
	function automatic hpdcache_pkg_is_amo_sc;
		// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_pkg.sv:137:40
		input reg [3:0] op;
		// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_pkg.sv:138:9
		case (op)
			4'h5: hpdcache_pkg_is_amo_sc = 1'b1;
			default: hpdcache_pkg_is_amo_sc = 1'b0;
		endcase
	endfunction
	assign st1_req_is_amo_sc = hpdcache_pkg_is_amo_sc(st1_req[4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))-:((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) >= ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) ? ((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) + 1 : (((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) - (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) + 1)]);
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:376:5
	function automatic hpdcache_pkg_is_amo_swap;
		// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_pkg.sv:144:42
		input reg [3:0] op;
		// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_pkg.sv:145:9
		case (op)
			4'h6: hpdcache_pkg_is_amo_swap = 1'b1;
			default: hpdcache_pkg_is_amo_swap = 1'b0;
		endcase
	endfunction
	assign st1_req_is_amo_swap = hpdcache_pkg_is_amo_swap(st1_req[4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))-:((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) >= ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) ? ((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) + 1 : (((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) - (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) + 1)]);
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:377:5
	function automatic hpdcache_pkg_is_amo_add;
		// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_pkg.sv:151:41
		input reg [3:0] op;
		// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_pkg.sv:152:9
		case (op)
			4'h7: hpdcache_pkg_is_amo_add = 1'b1;
			default: hpdcache_pkg_is_amo_add = 1'b0;
		endcase
	endfunction
	assign st1_req_is_amo_add = hpdcache_pkg_is_amo_add(st1_req[4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))-:((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) >= ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) ? ((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) + 1 : (((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) - (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) + 1)]);
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:378:5
	function automatic hpdcache_pkg_is_amo_and;
		// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_pkg.sv:158:41
		input reg [3:0] op;
		// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_pkg.sv:159:9
		case (op)
			4'h8: hpdcache_pkg_is_amo_and = 1'b1;
			default: hpdcache_pkg_is_amo_and = 1'b0;
		endcase
	endfunction
	assign st1_req_is_amo_and = hpdcache_pkg_is_amo_and(st1_req[4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))-:((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) >= ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) ? ((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) + 1 : (((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) - (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) + 1)]);
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:379:5
	function automatic hpdcache_pkg_is_amo_or;
		// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_pkg.sv:165:40
		input reg [3:0] op;
		// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_pkg.sv:166:9
		case (op)
			4'h9: hpdcache_pkg_is_amo_or = 1'b1;
			default: hpdcache_pkg_is_amo_or = 1'b0;
		endcase
	endfunction
	assign st1_req_is_amo_or = hpdcache_pkg_is_amo_or(st1_req[4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))-:((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) >= ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) ? ((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) + 1 : (((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) - (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) + 1)]);
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:380:5
	function automatic hpdcache_pkg_is_amo_xor;
		// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_pkg.sv:172:41
		input reg [3:0] op;
		// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_pkg.sv:173:9
		case (op)
			4'ha: hpdcache_pkg_is_amo_xor = 1'b1;
			default: hpdcache_pkg_is_amo_xor = 1'b0;
		endcase
	endfunction
	assign st1_req_is_amo_xor = hpdcache_pkg_is_amo_xor(st1_req[4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))-:((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) >= ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) ? ((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) + 1 : (((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) - (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) + 1)]);
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:381:5
	function automatic hpdcache_pkg_is_amo_max;
		// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_pkg.sv:179:41
		input reg [3:0] op;
		// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_pkg.sv:180:9
		case (op)
			4'hb: hpdcache_pkg_is_amo_max = 1'b1;
			default: hpdcache_pkg_is_amo_max = 1'b0;
		endcase
	endfunction
	assign st1_req_is_amo_max = hpdcache_pkg_is_amo_max(st1_req[4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))-:((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) >= ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) ? ((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) + 1 : (((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) - (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) + 1)]);
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:382:5
	function automatic hpdcache_pkg_is_amo_maxu;
		// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_pkg.sv:186:42
		input reg [3:0] op;
		// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_pkg.sv:187:9
		case (op)
			4'hc: hpdcache_pkg_is_amo_maxu = 1'b1;
			default: hpdcache_pkg_is_amo_maxu = 1'b0;
		endcase
	endfunction
	assign st1_req_is_amo_maxu = hpdcache_pkg_is_amo_maxu(st1_req[4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))-:((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) >= ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) ? ((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) + 1 : (((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) - (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) + 1)]);
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:383:5
	function automatic hpdcache_pkg_is_amo_min;
		// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_pkg.sv:193:41
		input reg [3:0] op;
		// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_pkg.sv:194:9
		case (op)
			4'hd: hpdcache_pkg_is_amo_min = 1'b1;
			default: hpdcache_pkg_is_amo_min = 1'b0;
		endcase
	endfunction
	assign st1_req_is_amo_min = hpdcache_pkg_is_amo_min(st1_req[4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))-:((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) >= ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) ? ((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) + 1 : (((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) - (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) + 1)]);
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:384:5
	function automatic hpdcache_pkg_is_amo_minu;
		// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_pkg.sv:200:42
		input reg [3:0] op;
		// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_pkg.sv:201:9
		case (op)
			4'he: hpdcache_pkg_is_amo_minu = 1'b1;
			default: hpdcache_pkg_is_amo_minu = 1'b0;
		endcase
	endfunction
	assign st1_req_is_amo_minu = hpdcache_pkg_is_amo_minu(st1_req[4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))-:((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) >= ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) ? ((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) + 1 : (((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) - (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) + 1)]);
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:385:5
	assign st1_req_is_cmo_inval = hpdcache_pkg_is_cmo_inval(st1_req[4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))-:((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) >= ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) ? ((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) + 1 : (((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) - (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) + 1)], st1_req[3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))-:((3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) >= (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) ? ((3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))) + 1 : ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) - (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) + 1)]);
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:386:5
	assign st1_req_is_cmo_fence = hpdcache_pkg_is_cmo_fence(st1_req[4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))-:((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) >= ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) ? ((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) + 1 : (((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) - (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) + 1)], st1_req[3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))-:((3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) >= (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) ? ((3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))) + 1 : ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) - (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) + 1)]);
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:387:5
	assign st1_req_is_cmo_prefetch = hpdcache_pkg_is_cmo_prefetch(st1_req[4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))-:((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) >= ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) ? ((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) + 1 : (((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) - (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) + 1)], st1_req[3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))-:((3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) >= (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) ? ((3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))) + 1 : ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) - (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) + 1)]);
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:392:5
	hpdcache_ctrl_pe hpdcache_ctrl_pe_i(
		.core_req_valid_i(core_req_valid_i),
		.core_req_ready_o(core_req_ready_o),
		.rtab_req_valid_i(st0_rtab_pop_try_valid),
		.rtab_req_ready_o(st0_rtab_pop_try_ready),
		.refill_req_valid_i(refill_req_valid_i),
		.refill_req_ready_o(refill_req_ready_o),
		.st0_req_is_uncacheable_i(st0_req_is_uncacheable),
		.st0_req_need_rsp_i(st0_req[2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)]),
		.st0_req_is_load_i(st0_req_is_load),
		.st0_req_is_store_i(st0_req_is_store),
		.st0_req_is_amo_i(st0_req_is_amo),
		.st0_req_is_cmo_fence_i(st0_req_is_cmo_fence),
		.st0_req_is_cmo_inval_i(st0_req_is_cmo_inval),
		.st0_req_is_cmo_prefetch_i(st0_req_is_cmo_prefetch),
		.st0_req_mshr_check_o(miss_mshr_check_o),
		.st0_req_cachedir_read_o(st0_req_cachedir_read),
		.st0_req_cachedata_read_o(st0_req_cachedata_read),
		.st1_req_valid_i(st1_req_valid_q),
		.st1_req_abort_i(st1_req_abort),
		.st1_req_rtab_i(st1_req_rtab_q),
		.st1_req_is_uncacheable_i(st1_req_is_uncacheable),
		.st1_req_need_rsp_i(st1_req[2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)]),
		.st1_req_is_load_i(st1_req_is_load),
		.st1_req_is_store_i(st1_req_is_store),
		.st1_req_is_amo_i(st1_req_is_amo),
		.st1_req_is_cmo_inval_i(st1_req_is_cmo_inval),
		.st1_req_is_cmo_fence_i(st1_req_is_cmo_fence),
		.st1_req_is_cmo_prefetch_i(st1_req_is_cmo_prefetch),
		.st1_req_valid_o(st1_req_valid_d),
		.st1_rsp_valid_o(st1_rsp_valid),
		.st1_rsp_aborted_o(st1_rsp_aborted),
		.st1_req_cachedir_updt_lru_o(st1_req_updt_lru),
		.st1_req_cachedata_write_o(st1_req_cachedata_write),
		.st1_req_cachedata_write_enable_o(st1_req_cachedata_write_enable),
		.st2_req_valid_i(st2_req_valid_q),
		.st2_req_is_prefetch_i(st2_req_is_prefetch_q),
		.st2_req_valid_o(st2_req_valid_d),
		.st2_req_we_o(st2_req_we),
		.st2_req_is_prefetch_o(st2_req_is_prefetch_d),
		.st2_req_mshr_alloc_o(miss_mshr_alloc_o),
		.st2_req_mshr_alloc_cs_o(miss_mshr_alloc_cs_o),
		.rtab_full_i(rtab_full),
		.rtab_check_o(st1_rtab_check),
		.rtab_check_hit_i(st1_rtab_check_hit),
		.st1_rtab_alloc_o(st1_rtab_alloc),
		.st1_rtab_alloc_and_link_o(st1_rtab_alloc_and_link),
		.st1_rtab_commit_o(st1_rtab_pop_try_commit),
		.st1_rtab_rback_o(st1_rtab_pop_try_rback),
		.st1_rtab_mshr_hit_o(st1_rtab_mshr_hit),
		.st1_rtab_mshr_full_o(st1_rtab_mshr_full),
		.st1_rtab_mshr_ready_o(st1_rtab_mshr_ready),
		.st1_rtab_wbuf_hit_o(st1_rtab_wbuf_hit),
		.st1_rtab_wbuf_not_ready_o(st1_rtab_wbuf_not_ready),
		.cachedir_hit_i(cachedir_hit_o),
		.cachedir_init_ready_i(hpdcache_init_ready),
		.mshr_alloc_ready_i(miss_mshr_alloc_ready_i),
		.mshr_hit_i(miss_mshr_hit_i),
		.mshr_full_i(miss_mshr_alloc_full_i),
		.refill_busy_i(refill_busy_i),
		.refill_core_rsp_valid_i(refill_core_rsp_valid_i),
		.wbuf_write_valid_o(wbuf_write_o),
		.wbuf_write_ready_i(wbuf_write_ready_i),
		.wbuf_read_hit_i(wbuf_read_hit_i),
		.wbuf_write_uncacheable_o(wbuf_write_uncacheable_o),
		.wbuf_read_flush_hit_o(wbuf_read_flush_hit_o),
		.uc_busy_i(uc_busy_i),
		.uc_req_valid_o(uc_req_valid_o),
		.uc_core_rsp_ready_o(uc_core_rsp_ready_o),
		.cmo_busy_i(cmo_busy_i),
		.cmo_wait_i(cmo_wait_i),
		.cmo_req_valid_o(cmo_req_valid_o),
		.evt_cache_write_miss_o(evt_cache_write_miss_o),
		.evt_cache_read_miss_o(evt_cache_read_miss_o),
		.evt_uncached_req_o(evt_uncached_req_o),
		.evt_cmo_req_o(evt_cmo_req_o),
		.evt_write_req_o(evt_write_req_o),
		.evt_read_req_o(evt_read_req_o),
		.evt_prefetch_req_o(evt_prefetch_req_o),
		.evt_req_on_hold_o(evt_req_on_hold_o),
		.evt_rtab_rollback_o(evt_rtab_rollback_o),
		.evt_stall_refill_o(evt_stall_refill_o),
		.evt_stall_o(evt_stall_o)
	);
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:489:5
	assign ctrl_empty_o = ~(st1_req_valid_q | st2_req_valid_q);
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:495:5
	localparam integer hpdcache_rtab_i_sv2v_pfunc_EB1A5 = $clog2($signed(HPDcacheCfg[671-:32]));
	hpdcache_rtab_6946D_40145 #(
		.hpdcache_nline_t_hpdcache_nline_t_HPDcacheCfg(hpdcache_nline_t_HPDcacheCfg),
		.hpdcache_req_addr_t_hpdcache_req_addr_t_HPDcacheCfg(hpdcache_req_addr_t_HPDcacheCfg),
		.rtab_entry_t_hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg(hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg),
		.rtab_ptr_t_hpdcache_rtab_i_sv2v_pfunc_EB1A5(hpdcache_rtab_i_sv2v_pfunc_EB1A5),
		.HPDcacheCfg(HPDcacheCfg)
	) hpdcache_rtab_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.empty_o(rtab_empty_o),
		.full_o(rtab_full),
		.check_i(st1_rtab_check),
		.check_nline_i(st1_req_nline),
		.check_hit_o(st1_rtab_check_hit),
		.alloc_i(st1_rtab_alloc),
		.alloc_and_link_i(st1_rtab_alloc_and_link),
		.alloc_req_i(st1_req),
		.alloc_mshr_hit_i(st1_rtab_mshr_hit),
		.alloc_mshr_full_i(st1_rtab_mshr_full),
		.alloc_mshr_ready_i(st1_rtab_mshr_ready),
		.alloc_wbuf_hit_i(st1_rtab_wbuf_hit),
		.alloc_wbuf_not_ready_i(st1_rtab_wbuf_not_ready),
		.pop_try_valid_o(st0_rtab_pop_try_valid),
		.pop_try_i(st0_rtab_pop_try_ready),
		.pop_try_req_o(st0_rtab_pop_try_req),
		.pop_try_ptr_o(st0_rtab_pop_try_ptr),
		.pop_commit_i(st1_rtab_pop_try_commit),
		.pop_commit_ptr_i(st1_rtab_pop_try_ptr_q),
		.pop_rback_i(st1_rtab_pop_try_rback),
		.pop_rback_ptr_i(st1_rtab_pop_try_ptr_q),
		.pop_rback_mshr_hit_i(st1_rtab_mshr_hit),
		.pop_rback_mshr_full_i(st1_rtab_mshr_full),
		.pop_rback_mshr_ready_i(st1_rtab_mshr_ready),
		.pop_rback_wbuf_hit_i(st1_rtab_wbuf_hit),
		.pop_rback_wbuf_not_ready_i(st1_rtab_wbuf_not_ready),
		.wbuf_addr_o(wbuf_rtab_addr_o),
		.wbuf_is_read_o(wbuf_rtab_is_read_o),
		.wbuf_hit_open_i(wbuf_rtab_hit_open_i),
		.wbuf_hit_pend_i(wbuf_rtab_hit_pend_i),
		.wbuf_hit_sent_i(wbuf_rtab_hit_sent_i),
		.wbuf_not_ready_i(wbuf_rtab_not_ready_i),
		.miss_ready_i(miss_mshr_alloc_ready_i),
		.refill_i(refill_updt_rtab_i),
		.refill_nline_i(refill_nline_i),
		.cfg_single_entry_i(cfg_rtab_single_entry_i)
	);
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:555:5
	always @(posedge clk_i) begin : st1_req_payload_ff
		// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:557:9
		if (core_req_ready_o | st0_rtab_pop_try_ready)
			// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:558:13
			st1_req_q <= st0_req;
	end
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:562:5
	always @(posedge clk_i or negedge rst_ni) begin : st1_req_valid_ff
		// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:564:9
		if (!rst_ni) begin
			// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:565:13
			st1_req_valid_q <= 1'b0;
			// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:566:13
			st1_req_rtab_q <= 1'b0;
			// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:567:13
			st1_rtab_pop_try_ptr_q <= 1'sb0;
		end
		else begin
			// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:570:13
			st1_req_valid_q <= st1_req_valid_d;
			// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:571:13
			if (core_req_ready_o | st0_rtab_pop_try_ready) begin
				// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:572:17
				st1_req_rtab_q <= st0_rtab_pop_try_ready;
				// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:573:17
				if (st0_rtab_pop_try_ready)
					// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:574:21
					st1_rtab_pop_try_ptr_q <= st0_rtab_pop_try_ptr;
			end
		end
	end
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:583:5
	always @(posedge clk_i) begin : st2_req_payload_ff
		// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:585:9
		if (st2_req_we) begin
			// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:586:13
			st2_req_need_rsp_q <= st1_req[2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)];
			// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:587:13
			st2_req_addr_q <= st1_req_addr;
			// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:588:13
			st2_req_sid_q <= st1_req[hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))-:((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))) >= (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))) ? ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))) - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) + 1 : ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))) - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) + 1)];
			// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:589:13
			st2_req_tid_q <= st1_req[hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))-:((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))) >= (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)) ? ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))) - (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))) + 1 : ((2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)) - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))) + 1)];
		end
	end
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:593:5
	always @(posedge clk_i or negedge rst_ni) begin : st2_req_valid_ff
		// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:595:9
		if (!rst_ni) begin
			// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:596:13
			st2_req_valid_q <= 1'b0;
			// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:597:13
			st2_req_is_prefetch_q <= 1'b0;
		end
		else begin
			// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:599:13
			st2_req_valid_q <= st2_req_valid_d;
			// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:600:13
			st2_req_is_prefetch_q <= st2_req_is_prefetch_d;
		end
	end
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:607:5
	assign st0_req_set = st0_req[(hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] - 1) - HPDcacheCfg[447-:32])+:HPDcacheCfg[415-:32]];
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:608:5
	assign st0_req_word = st0_req[(hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] - 1) - HPDcacheCfg[479-:32])+:HPDcacheCfg[511-:32]];
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:611:5
	assign st1_req_set = st1_req[(hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] - 1) - HPDcacheCfg[447-:32])+:HPDcacheCfg[415-:32]];
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:612:5
	assign st1_req_word = st1_req[(hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] - 1) - HPDcacheCfg[479-:32])+:HPDcacheCfg[511-:32]];
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:614:5
	assign st1_req_addr = {st1_req[hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1-:((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1) >= 2 ? hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 0 : 3 - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))], st1_req[hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))-:((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))) >= ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))))) ? ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))))) + 1 : (((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))))) - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))))) + 1)]};
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:615:5
	assign st1_req_nline = st1_req_addr[HPDcacheCfg[447-:32]+:HPDcacheCfg[383-:32]];
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:617:5
	assign st2_req_word = st2_req_addr_q[HPDcacheCfg[479-:32]+:HPDcacheCfg[511-:32]];
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:620:5
	hpdcache_memctrl_712A3_4BE95 #(
		.hpdcache_data_be_t_hpdcache_data_be_t_hpdcache_data_be_t_hpdcache_data_be_t_HPDcacheCfg(hpdcache_data_be_t_hpdcache_data_be_t_hpdcache_data_be_t_HPDcacheCfg),
		.hpdcache_data_word_t_hpdcache_data_word_t_hpdcache_data_word_t_hpdcache_data_word_t_HPDcacheCfg(hpdcache_data_word_t_hpdcache_data_word_t_hpdcache_data_word_t_HPDcacheCfg),
		.hpdcache_dir_entry_t_hpdcache_dir_entry_t_hpdcache_tag_t_hpdcache_tag_t_HPDcacheCfg(hpdcache_dir_entry_t_hpdcache_tag_t_hpdcache_tag_t_HPDcacheCfg),
		.hpdcache_nline_t_hpdcache_nline_t_HPDcacheCfg(hpdcache_nline_t_HPDcacheCfg),
		.hpdcache_refill_be_t_hpdcache_refill_be_t_HPDcacheCfg(hpdcache_refill_be_t_HPDcacheCfg),
		.hpdcache_refill_be_t_hpdcache_refill_be_t_hpdcache_data_be_t_hpdcache_data_be_t_HPDcacheCfg(hpdcache_refill_be_t_hpdcache_data_be_t_hpdcache_data_be_t_HPDcacheCfg),
		.hpdcache_refill_data_t_hpdcache_refill_data_t_HPDcacheCfg(hpdcache_refill_data_t_HPDcacheCfg),
		.hpdcache_refill_data_t_hpdcache_refill_data_t_hpdcache_data_word_t_hpdcache_data_word_t_HPDcacheCfg(hpdcache_refill_data_t_hpdcache_data_word_t_hpdcache_data_word_t_HPDcacheCfg),
		.hpdcache_req_be_t_hpdcache_req_be_t_hpdcache_req_be_t_hpdcache_req_be_t_HPDcacheCfg(hpdcache_req_be_t_hpdcache_req_be_t_hpdcache_req_be_t_HPDcacheCfg),
		.hpdcache_req_data_t_hpdcache_req_data_t_hpdcache_req_data_t_hpdcache_req_data_t_HPDcacheCfg(hpdcache_req_data_t_hpdcache_req_data_t_hpdcache_req_data_t_HPDcacheCfg),
		.hpdcache_set_t_hpdcache_set_t_HPDcacheCfg(hpdcache_set_t_HPDcacheCfg),
		.hpdcache_tag_t_hpdcache_tag_t_hpdcache_tag_t_hpdcache_tag_t_HPDcacheCfg(hpdcache_tag_t_hpdcache_tag_t_hpdcache_tag_t_HPDcacheCfg),
		.hpdcache_way_vector_t_hpdcache_way_vector_t_HPDcacheCfg(hpdcache_way_vector_t_HPDcacheCfg),
		.hpdcache_word_t_hpdcache_word_t_HPDcacheCfg(hpdcache_word_t_HPDcacheCfg),
		.HPDcacheCfg(HPDcacheCfg)
	) hpdcache_memctrl_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.ready_o(hpdcache_init_ready),
		.dir_match_i(st0_req_cachedir_read),
		.dir_match_set_i(st0_req_set),
		.dir_match_tag_i(st1_req[hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1-:((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1) >= 2 ? hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 0 : 3 - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))]),
		.dir_update_lru_i(st1_req_updt_lru),
		.dir_hit_way_o(st1_dir_hit),
		.dir_amo_match_i(uc_dir_amo_match_i),
		.dir_amo_match_set_i(uc_dir_amo_match_set_i),
		.dir_amo_match_tag_i(uc_dir_amo_match_tag_i),
		.dir_amo_update_plru_i(uc_dir_amo_update_plru_i),
		.dir_amo_hit_way_o(uc_dir_amo_hit_way_o),
		.dir_refill_sel_victim_i(refill_sel_victim_i),
		.dir_refill_i(refill_write_dir_i),
		.dir_refill_set_i(refill_set_i),
		.dir_refill_entry_i(refill_dir_entry_i),
		.dir_refill_updt_plru_i(refill_updt_plru_i),
		.dir_victim_way_o(refill_victim_way_o),
		.dir_inval_check_i(inval_check_dir_i),
		.dir_inval_nline_i(inval_nline_i),
		.dir_inval_write_i(inval_write_dir_i),
		.dir_inval_hit_o(inval_hit_o),
		.dir_cmo_check_i(cmo_dir_check_i),
		.dir_cmo_check_set_i(cmo_dir_check_set_i),
		.dir_cmo_check_tag_i(cmo_dir_check_tag_i),
		.dir_cmo_check_hit_way_o(cmo_dir_check_hit_way_o),
		.dir_cmo_inval_i(cmo_dir_inval_i),
		.dir_cmo_inval_set_i(cmo_dir_inval_set_i),
		.dir_cmo_inval_way_i(cmo_dir_inval_way_i),
		.data_req_read_i(st0_req_cachedata_read),
		.data_req_read_set_i(st0_req_set),
		.data_req_read_size_i(st0_req[3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))-:((3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) >= (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) ? ((3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))) + 1 : ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) - (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) + 1)]),
		.data_req_read_word_i(st0_req_word),
		.data_req_read_data_o(st1_read_data),
		.data_req_write_i(st1_req_cachedata_write),
		.data_req_write_enable_i(st1_req_cachedata_write_enable),
		.data_req_write_set_i(st1_req_set),
		.data_req_write_size_i(st1_req[3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))-:((3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) >= (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) ? ((3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))) + 1 : ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) - (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) + 1)]),
		.data_req_write_word_i(st1_req_word),
		.data_req_write_data_i(st1_req[(hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))-:(((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) >= (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) ? (((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) - (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))))) + 1 : ((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))) + 1)]),
		.data_req_write_be_i(st1_req[(hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))-:(((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) >= (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))) ? (((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) - (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) + 1 : ((3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) + 1)]),
		.data_amo_write_i(uc_data_amo_write_i),
		.data_amo_write_enable_i(uc_data_amo_write_enable_i),
		.data_amo_write_set_i(uc_data_amo_write_set_i),
		.data_amo_write_size_i(uc_data_amo_write_size_i),
		.data_amo_write_word_i(uc_data_amo_write_word_i),
		.data_amo_write_data_i(uc_data_amo_write_data_i),
		.data_amo_write_be_i(uc_data_amo_write_be_i),
		.data_refill_i(refill_write_data_i),
		.data_refill_way_i(refill_victim_way_i),
		.data_refill_set_i(refill_set_i),
		.data_refill_word_i(refill_word_i),
		.data_refill_data_i(refill_data_i)
	);
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:702:5
	assign cachedir_hit_o = |st1_dir_hit;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:707:5
	assign wbuf_write_addr_o = st1_req_addr;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:708:5
	assign wbuf_write_data_o = st1_req[(hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))-:(((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) >= (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) ? (((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) - (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))))) + 1 : ((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))) + 1)];
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:709:5
	assign wbuf_write_be_o = st1_req[(hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))-:(((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) >= (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))) ? (((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) - (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) + 1 : ((3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) + 1)];
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:710:5
	assign wbuf_flush_all_o = (cmo_wbuf_flush_all_i | uc_wbuf_flush_all_i) | wbuf_flush_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:715:5
	assign miss_mshr_check_offset_o = st0_req[hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))-:((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))) >= ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))))) ? ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))))) + 1 : (((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))))) - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))))) + 1)];
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:716:5
	assign miss_mshr_check_nline_o = st1_req_nline;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:717:5
	assign miss_mshr_alloc_nline_o = st2_req_addr_q[HPDcacheCfg[447-:32]+:HPDcacheCfg[383-:32]];
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:719:5
	assign miss_mshr_alloc_tid_o = st2_req_tid_q;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:720:5
	assign miss_mshr_alloc_sid_o = st2_req_sid_q;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:721:5
	assign miss_mshr_alloc_word_o = st2_req_word;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:722:5
	assign miss_mshr_alloc_need_rsp_o = st2_req_need_rsp_q;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:723:5
	assign miss_mshr_alloc_is_prefetch_o = st2_req_is_prefetch_q;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:728:5
	assign uc_lrsc_snoop_o = st1_req_valid_q & st1_req_is_store;
	assign uc_lrsc_snoop_addr_o = st1_req_addr;
	assign uc_lrsc_snoop_size_o = st1_req[3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))-:((3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) >= (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) ? ((3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))) + 1 : ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) - (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) + 1)];
	assign uc_req_addr_o = st1_req_addr;
	assign uc_req_size_o = st1_req[3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))-:((3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) >= (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) ? ((3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))) + 1 : ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) - (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) + 1)];
	assign uc_req_data_o = st1_req[(hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))-:(((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) >= (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) ? (((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) - (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))))) + 1 : ((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))) + 1)];
	assign uc_req_be_o = st1_req[(hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))-:(((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) >= (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))) ? (((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) - (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) + 1 : ((3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) + 1)];
	assign uc_req_uc_o = st1_req_is_uncacheable;
	assign uc_req_sid_o = st1_req[hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))-:((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))) >= (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))) ? ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))) - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) + 1 : ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))) - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) + 1)];
	assign uc_req_tid_o = st1_req[hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))-:((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))) >= (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)) ? ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))) - (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))) + 1 : ((2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)) - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))) + 1)];
	assign uc_req_need_rsp_o = st1_req[2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)];
	assign uc_req_op_o[12] = st1_req_is_load;
	assign uc_req_op_o[11] = st1_req_is_store;
	assign uc_req_op_o[10] = st1_req_is_amo_lr;
	assign uc_req_op_o[9] = st1_req_is_amo_sc;
	assign uc_req_op_o[8] = st1_req_is_amo_swap;
	assign uc_req_op_o[7] = st1_req_is_amo_add;
	assign uc_req_op_o[6] = st1_req_is_amo_and;
	assign uc_req_op_o[5] = st1_req_is_amo_or;
	assign uc_req_op_o[4] = st1_req_is_amo_xor;
	assign uc_req_op_o[3] = st1_req_is_amo_max;
	assign uc_req_op_o[2] = st1_req_is_amo_maxu;
	assign uc_req_op_o[1] = st1_req_is_amo_min;
	assign uc_req_op_o[0] = st1_req_is_amo_minu;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:756:5
	assign cmo_req_addr_o = st1_req_addr;
	assign cmo_req_wdata_o = st1_req[(hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))-:(((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) >= (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) ? (((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) - (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))))) + 1 : ((4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) - ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))) + 1)];
	assign cmo_req_op_o[0] = st1_req_is_cmo_fence;
	function automatic hpdcache_pkg_is_cmo_inval_by_nline;
		// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_pkg.sv:228:52
		input reg [2:0] sz;
		// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_pkg.sv:229:9
		hpdcache_pkg_is_cmo_inval_by_nline = sz == 3'h2;
	endfunction
	assign cmo_req_op_o[3] = st1_req_is_cmo_inval & hpdcache_pkg_is_cmo_inval_by_nline(st1_req[3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))-:((3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) >= (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) ? ((3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))) + 1 : ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) - (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) + 1)]);
	function automatic hpdcache_pkg_is_cmo_inval_by_set;
		// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_pkg.sv:232:50
		input reg [2:0] sz;
		// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_pkg.sv:233:9
		hpdcache_pkg_is_cmo_inval_by_set = sz == 3'h3;
	endfunction
	assign cmo_req_op_o[2] = st1_req_is_cmo_inval & hpdcache_pkg_is_cmo_inval_by_set(st1_req[3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))-:((3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) >= (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) ? ((3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))) + 1 : ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) - (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) + 1)]);
	function automatic hpdcache_pkg_is_cmo_inval_all;
		// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_pkg.sv:236:47
		input reg [2:0] sz;
		// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_pkg.sv:237:9
		hpdcache_pkg_is_cmo_inval_all = sz == 3'h4;
	endfunction
	assign cmo_req_op_o[1] = st1_req_is_cmo_inval & hpdcache_pkg_is_cmo_inval_all(st1_req[3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))-:((3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) >= (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) ? ((3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))) + 1 : ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) - (3 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) + 1)]);
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:769:5
	assign core_rsp_valid_o = (refill_core_rsp_valid_i | (uc_core_rsp_valid_i & uc_core_rsp_ready_o)) | st1_rsp_valid;
	assign core_rsp_o[(hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1157-:32] * hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1285-:32]) + (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32] + (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1))-:(((hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1157-:32] * hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1285-:32]) + (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32] + (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1))) >= (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32] + (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 2)) ? (((hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1157-:32] * hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1285-:32]) + (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32] + (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1))) - (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32] + (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 2))) + 1 : ((hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32] + (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 2)) - ((hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1157-:32] * hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1285-:32]) + (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32] + (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1)))) + 1)] = (refill_core_rsp_valid_i ? refill_core_rsp_i[(hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1157-:32] * hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1285-:32]) + (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32] + (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1))-:(((hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1157-:32] * hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1285-:32]) + (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32] + (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1))) >= (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32] + (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 2)) ? (((hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1157-:32] * hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1285-:32]) + (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32] + (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1))) - (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32] + (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 2))) + 1 : ((hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32] + (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 2)) - ((hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1157-:32] * hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1285-:32]) + (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32] + (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1)))) + 1)] : (uc_core_rsp_valid_i ? uc_core_rsp_i[(hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1157-:32] * hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1285-:32]) + (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32] + (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1))-:(((hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1157-:32] * hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1285-:32]) + (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32] + (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1))) >= (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32] + (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 2)) ? (((hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1157-:32] * hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1285-:32]) + (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32] + (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1))) - (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32] + (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 2))) + 1 : ((hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32] + (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 2)) - ((hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1157-:32] * hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1285-:32]) + (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32] + (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1)))) + 1)] : st1_read_data));
	assign core_rsp_o[hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32] + (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1)-:((hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32] + (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1)) >= (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 2) ? ((hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32] + (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1)) - (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 2)) + 1 : ((hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 2) - (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32] + (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1))) + 1)] = (refill_core_rsp_valid_i ? refill_core_rsp_i[hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32] + (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1)-:((hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32] + (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1)) >= (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 2) ? ((hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32] + (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1)) - (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 2)) + 1 : ((hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 2) - (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32] + (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1))) + 1)] : (uc_core_rsp_valid_i ? uc_core_rsp_i[hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32] + (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1)-:((hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32] + (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1)) >= (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 2) ? ((hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32] + (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1)) - (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 2)) + 1 : ((hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 2) - (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32] + (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1))) + 1)] : st1_req[hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))-:((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))) >= (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))) ? ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))) - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) + 1 : ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))) - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) + 1)]));
	assign core_rsp_o[hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1-:((hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1) >= 2 ? hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 0 : 3 - (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1))] = (refill_core_rsp_valid_i ? refill_core_rsp_i[hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1-:((hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1) >= 2 ? hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 0 : 3 - (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1))] : (uc_core_rsp_valid_i ? uc_core_rsp_i[hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1-:((hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1) >= 2 ? hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 0 : 3 - (hpdcache_rsp_t_hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1))] : st1_req[hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))-:((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))) >= (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)) ? ((hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))) - (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))) + 1 : ((2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)) - (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))) + 1)]));
	assign core_rsp_o[1] = (refill_core_rsp_valid_i ? refill_core_rsp_i[1] : (uc_core_rsp_valid_i ? uc_core_rsp_i[1] : 1'b0));
	assign core_rsp_o[0] = st1_rsp_aborted;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:790:5
	// removed an assertion item
	// assert property (@(posedge clk_i) disable iff (!rst_ni)
	// 	$onehot0({core_req_ready_o, st0_rtab_pop_try_ready, refill_req_ready_o})
	// ) else begin
	// 	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:792:21
	// 	$error("ctrl: only one request can be served per cycle");
	// end
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:794:5
	// removed an assertion item
	// property prop_core_req_size_max;
	// 	@(posedge clk_i) disable iff (!rst_ni)
	// 		((core_req_valid_i && core_req_ready_o) && (core_req_i.op != hpdcache_pkg_HPDCACHE_REQ_CMO) |-> (2 ** core_req_i.size) <= HPDcacheCfg.reqDataBytes)
	// endproperty
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:803:5
	// removed an assertion item
	// assert property (
	// 	prop_core_req_size_max
	// ) else begin
	// 	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:804:13
	// 	$error("ctrl: bad SIZE for request");
	// end
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:806:5
	function automatic signed [31:0] sv2v_cast_32_signed;
		input reg signed [31:0] inp;
		sv2v_cast_32_signed = inp;
	endfunction
	function automatic check_is_be_aligned;
		// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:807:7
		input reg [hpdcache_req_offset_t_hpdcache_req_offset_t_hpdcache_req_offset_t_HPDcacheCfg[287-:32] - 1:0] req_offset;
		// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:808:7
		input reg [(hpdcache_req_be_t_hpdcache_req_be_t_hpdcache_req_be_t_HPDcacheCfg[1157-:32] * (hpdcache_req_be_t_hpdcache_req_be_t_hpdcache_req_be_t_HPDcacheCfg[1285-:32] / 8)) - 1:0] req_be;
		// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:810:9
		reg signed [31:0] offset;
		begin
			offset = sv2v_cast_32_signed(req_offset) % HPDcacheCfg[223-:32];
			// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:811:9
			check_is_be_aligned = ((req_be >> offset) << offset) == req_be;
		end
	endfunction
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:814:5
	// removed an assertion item
	// property prop_core_req_be_align;
	// 	@(posedge clk_i) disable iff (!rst_ni)
	// 		((core_req_valid_i && core_req_ready_o) && (hpdcache_pkg_is_store(core_req_i.op) || hpdcache_pkg_is_amo(core_req_i.op)) |-> check_is_be_aligned(core_req_i.addr_offset, core_req_i.be))
	// endproperty
	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:823:5
	// removed an assertion item
	// assert property (
	// 	prop_core_req_be_align
	// ) else begin
	// 	// Trace: core/cache_subsystem/hpdcache/rtl/src/hpdcache_ctrl.sv:824:13
	// 	$error("ctrl: bad BE alignment for request");
	// end
endmodule
