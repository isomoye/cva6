module frontend_FEAA5_C53EA (
	clk_i,
	rst_ni,
	boot_addr_i,
	flush_bp_i,
	flush_i,
	halt_i,
	set_pc_commit_i,
	pc_commit_i,
	ex_valid_i,
	resolved_branch_i,
	eret_i,
	epc_i,
	trap_vector_base_i,
	set_debug_pc_i,
	debug_mode_i,
	icache_dreq_o,
	icache_dreq_i,
	fetch_entry_o,
	fetch_entry_valid_o,
	fetch_entry_ready_i
);
	// removed localparam type bp_resolve_t_CVA6Cfg_type
	// removed localparam type bp_resolve_t_config_pkg_NrMaxRules_type
	parameter [17102:0] bp_resolve_t_CVA6Cfg = 0;
	parameter signed [31:0] bp_resolve_t_config_pkg_NrMaxRules = 0;
	// removed localparam type fetch_entry_t_CVA6Cfg_type
	// removed localparam type fetch_entry_t_config_pkg_NrMaxRules_type
	parameter [17102:0] fetch_entry_t_CVA6Cfg = 0;
	parameter signed [31:0] fetch_entry_t_config_pkg_NrMaxRules = 0;
	// removed localparam type icache_dreq_t_CVA6Cfg_type
	// removed localparam type icache_dreq_t_config_pkg_NrMaxRules_type
	parameter [17102:0] icache_dreq_t_CVA6Cfg = 0;
	parameter signed [31:0] icache_dreq_t_config_pkg_NrMaxRules = 0;
	// removed localparam type icache_drsp_t_CVA6Cfg_type
	// removed localparam type icache_drsp_t_config_pkg_NrMaxRules_type
	parameter [17102:0] icache_drsp_t_CVA6Cfg = 0;
	parameter signed [31:0] icache_drsp_t_config_pkg_NrMaxRules = 0;
	reg _sv2v_0;
	// removed import ariane_pkg::*;
	// Trace: core/frontend/frontend.sv:21:15
	localparam config_pkg_NrMaxRules = 16;
	// removed localparam type config_pkg_cache_type_t
	// removed localparam type config_pkg_noc_type_e
	// removed localparam type config_pkg_vm_mode_t
	// removed localparam type config_pkg_cva6_cfg_t
	localparam [17102:0] config_pkg_cva6_cfg_empty = 17103'd0;
	parameter [17102:0] CVA6Cfg = config_pkg_cva6_cfg_empty;
	// Trace: core/frontend/frontend.sv:22:20
	// removed localparam type bp_resolve_t
	// Trace: core/frontend/frontend.sv:23:20
	// removed localparam type fetch_entry_t
	// Trace: core/frontend/frontend.sv:24:20
	// removed localparam type icache_dreq_t
	// Trace: core/frontend/frontend.sv:25:20
	// removed localparam type icache_drsp_t
	// Trace: core/frontend/frontend.sv:28:5
	input wire clk_i;
	// Trace: core/frontend/frontend.sv:30:5
	input wire rst_ni;
	// Trace: core/frontend/frontend.sv:32:5
	input wire [CVA6Cfg[17070-:32] - 1:0] boot_addr_i;
	// Trace: core/frontend/frontend.sv:34:5
	input wire flush_bp_i;
	// Trace: core/frontend/frontend.sv:36:5
	input wire flush_i;
	// Trace: core/frontend/frontend.sv:38:5
	input wire halt_i;
	// Trace: core/frontend/frontend.sv:40:5
	input wire set_pc_commit_i;
	// Trace: core/frontend/frontend.sv:42:5
	input wire [CVA6Cfg[17070-:32] - 1:0] pc_commit_i;
	// Trace: core/frontend/frontend.sv:44:5
	input wire ex_valid_i;
	// Trace: core/frontend/frontend.sv:46:5
	input wire [((1 + bp_resolve_t_CVA6Cfg[9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + bp_resolve_t_CVA6Cfg[9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 4:0] resolved_branch_i;
	// Trace: core/frontend/frontend.sv:48:5
	input wire eret_i;
	// Trace: core/frontend/frontend.sv:50:5
	input wire [CVA6Cfg[17070-:32] - 1:0] epc_i;
	// Trace: core/frontend/frontend.sv:52:5
	input wire [CVA6Cfg[17070-:32] - 1:0] trap_vector_base_i;
	// Trace: core/frontend/frontend.sv:54:5
	input wire set_debug_pc_i;
	// Trace: core/frontend/frontend.sv:56:5
	input wire debug_mode_i;
	// Trace: core/frontend/frontend.sv:58:5
	output reg [(4 + icache_dreq_t_CVA6Cfg[9509 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) - 1:0] icache_dreq_o;
	// Trace: core/frontend/frontend.sv:60:5
	input wire [((((2 + icache_drsp_t_CVA6Cfg[643-:32]) + icache_drsp_t_CVA6Cfg[708-:32]) + icache_drsp_t_CVA6Cfg[9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + ((((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33) >= 0 ? ((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 34 : 1 - (((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33))) - 1:0] icache_dreq_i;
	// Trace: core/frontend/frontend.sv:62:5
	output wire [(CVA6Cfg[16841-:32] * (((fetch_entry_t_CVA6Cfg[9509 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 32) + (3 + fetch_entry_t_CVA6Cfg[9509 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)])) + ((((fetch_entry_t_CVA6Cfg[9541 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + fetch_entry_t_CVA6Cfg[9541 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + fetch_entry_t_CVA6Cfg[9445 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[9541 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + fetch_entry_t_CVA6Cfg[9541 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + fetch_entry_t_CVA6Cfg[9445 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[9541 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + fetch_entry_t_CVA6Cfg[9541 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + fetch_entry_t_CVA6Cfg[9445 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + (32 + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + ((fetch_entry_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33)))) - 1:0] fetch_entry_o;
	// Trace: core/frontend/frontend.sv:64:5
	output wire [CVA6Cfg[16841-:32] - 1:0] fetch_entry_valid_o;
	// Trace: core/frontend/frontend.sv:66:5
	input wire [CVA6Cfg[16841-:32] - 1:0] fetch_entry_ready_i;
	// Trace: core/frontend/frontend.sv:69:3
	// removed localparam type bht_update_t
	// Trace: core/frontend/frontend.sv:75:3
	// removed localparam type btb_prediction_t
	// Trace: core/frontend/frontend.sv:80:3
	// removed localparam type btb_update_t
	// Trace: core/frontend/frontend.sv:86:3
	// removed localparam type ras_t
	// Trace: core/frontend/frontend.sv:92:3
	reg [CVA6Cfg[643-:32] - 1:0] icache_data_q;
	// Trace: core/frontend/frontend.sv:93:3
	reg icache_valid_q;
	// Trace: core/frontend/frontend.sv:94:3
	// removed localparam type ariane_pkg_frontend_exception_t
	reg [1:0] icache_ex_valid_q;
	// Trace: core/frontend/frontend.sv:95:3
	reg [CVA6Cfg[17070-:32] - 1:0] icache_vaddr_q;
	// Trace: core/frontend/frontend.sv:96:3
	reg [CVA6Cfg[17006-:32] - 1:0] icache_gpaddr_q;
	// Trace: core/frontend/frontend.sv:97:3
	reg [31:0] icache_tinst_q;
	// Trace: core/frontend/frontend.sv:98:3
	reg icache_gva_q;
	// Trace: core/frontend/frontend.sv:99:3
	wire instr_queue_ready;
	// Trace: core/frontend/frontend.sv:100:3
	wire [CVA6Cfg[579-:32] - 1:0] instr_queue_consumed;
	// Trace: core/frontend/frontend.sv:102:3
	reg [(1 + CVA6Cfg[17070-:32]) - 1:0] btb_q;
	// Trace: core/frontend/frontend.sv:103:3
	// removed localparam type ariane_pkg_bht_prediction_t
	reg [1:0] bht_q;
	// Trace: core/frontend/frontend.sv:105:3
	wire if_ready;
	// Trace: core/frontend/frontend.sv:106:3
	reg [CVA6Cfg[17070-:32] - 1:0] npc_d;
	reg [CVA6Cfg[17070-:32] - 1:0] npc_q;
	// Trace: core/frontend/frontend.sv:109:3
	reg npc_rst_load_q;
	// Trace: core/frontend/frontend.sv:111:3
	wire replay;
	// Trace: core/frontend/frontend.sv:112:3
	wire [CVA6Cfg[17070-:32] - 1:0] replay_addr;
	// Trace: core/frontend/frontend.sv:115:3
	wire [$clog2(CVA6Cfg[579-:32]) - 1:0] shamt;
	// Trace: core/frontend/frontend.sv:117:3
	generate
		if (CVA6Cfg[16544]) begin : gen_shamt
			// Trace: core/frontend/frontend.sv:118:5
			assign shamt = icache_dreq_i[(icache_drsp_t_CVA6Cfg[9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (((((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33) >= 0 ? ((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 34 : 1 - (((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33)) - 1)) - ((icache_drsp_t_CVA6Cfg[9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1) - $clog2(CVA6Cfg[579-:32])):(icache_drsp_t_CVA6Cfg[9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (((((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33) >= 0 ? ((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 34 : 1 - (((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33)) - 1)) - (icache_drsp_t_CVA6Cfg[9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 2)];
		end
		else begin : genblk1
			// Trace: core/frontend/frontend.sv:120:5
			assign shamt = 1'b0;
		end
	endgenerate
	// Trace: core/frontend/frontend.sv:127:3
	wire [CVA6Cfg[579-:32] - 1:0] rvi_return;
	wire [CVA6Cfg[579-:32] - 1:0] rvi_call;
	wire [CVA6Cfg[579-:32] - 1:0] rvi_branch;
	wire [CVA6Cfg[579-:32] - 1:0] rvi_jalr;
	wire [CVA6Cfg[579-:32] - 1:0] rvi_jump;
	// Trace: core/frontend/frontend.sv:128:3
	wire [(CVA6Cfg[579-:32] * CVA6Cfg[17070-:32]) - 1:0] rvi_imm;
	// Trace: core/frontend/frontend.sv:130:3
	wire [CVA6Cfg[579-:32] - 1:0] rvc_branch;
	wire [CVA6Cfg[579-:32] - 1:0] rvc_jump;
	wire [CVA6Cfg[579-:32] - 1:0] rvc_jr;
	wire [CVA6Cfg[579-:32] - 1:0] rvc_return;
	wire [CVA6Cfg[579-:32] - 1:0] rvc_jalr;
	wire [CVA6Cfg[579-:32] - 1:0] rvc_call;
	// Trace: core/frontend/frontend.sv:131:3
	wire [(CVA6Cfg[579-:32] * CVA6Cfg[17070-:32]) - 1:0] rvc_imm;
	// Trace: core/frontend/frontend.sv:133:3
	wire [(CVA6Cfg[579-:32] * 32) - 1:0] instr;
	// Trace: core/frontend/frontend.sv:134:3
	wire [(CVA6Cfg[579-:32] * CVA6Cfg[17070-:32]) - 1:0] addr;
	// Trace: core/frontend/frontend.sv:135:3
	wire [CVA6Cfg[579-:32] - 1:0] instruction_valid;
	// Trace: core/frontend/frontend.sv:137:3
	wire [(CVA6Cfg[579-:32] * 2) - 1:0] bht_prediction;
	// Trace: core/frontend/frontend.sv:138:3
	wire [(CVA6Cfg[579-:32] * (1 + CVA6Cfg[17070-:32])) - 1:0] btb_prediction;
	// Trace: core/frontend/frontend.sv:139:3
	wire [(CVA6Cfg[579-:32] * 2) - 1:0] bht_prediction_shifted;
	// Trace: core/frontend/frontend.sv:140:3
	wire [(CVA6Cfg[579-:32] * (1 + CVA6Cfg[17070-:32])) - 1:0] btb_prediction_shifted;
	// Trace: core/frontend/frontend.sv:141:3
	wire [(1 + CVA6Cfg[17070-:32]) - 1:0] ras_predict;
	// Trace: core/frontend/frontend.sv:142:3
	wire [CVA6Cfg[17070-:32] - 1:0] vpc_btb;
	// Trace: core/frontend/frontend.sv:145:3
	wire is_mispredict;
	// Trace: core/frontend/frontend.sv:146:3
	reg ras_push;
	reg ras_pop;
	// Trace: core/frontend/frontend.sv:147:3
	reg [CVA6Cfg[17070-:32] - 1:0] ras_update;
	// Trace: core/frontend/frontend.sv:150:3
	reg [CVA6Cfg[17070-:32] - 1:0] predict_address;
	// Trace: core/frontend/frontend.sv:151:3
	// removed localparam type ariane_pkg_cf_t
	reg [(CVA6Cfg[579-:32] * 3) - 1:0] cf_type;
	// Trace: core/frontend/frontend.sv:152:3
	reg [CVA6Cfg[579-:32] - 1:0] taken_rvi_cf;
	// Trace: core/frontend/frontend.sv:153:3
	reg [CVA6Cfg[579-:32] - 1:0] taken_rvc_cf;
	// Trace: core/frontend/frontend.sv:155:3
	wire serving_unaligned;
	// Trace: core/frontend/frontend.sv:157:3
	instr_realign #(.CVA6Cfg(CVA6Cfg)) i_instr_realign(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(icache_dreq_o[icache_dreq_t_CVA6Cfg[9509 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 1]),
		.valid_i(icache_valid_q),
		.serving_unaligned_o(serving_unaligned),
		.address_i(icache_vaddr_q),
		.data_i(icache_data_q),
		.valid_o(instruction_valid),
		.addr_o(addr),
		.instr_o(instr)
	);
	// Trace: core/frontend/frontend.sv:177:3
	generate
		if (CVA6Cfg[16544]) begin : gen_btb_prediction_shifted
			// Trace: core/frontend/frontend.sv:178:5
			assign bht_prediction_shifted[0+:2] = (serving_unaligned ? bht_q : bht_prediction[addr[0 + ($clog2(CVA6Cfg[579-:32]) >= 1 ? $clog2(CVA6Cfg[579-:32]) : ($clog2(CVA6Cfg[579-:32]) + ($clog2(CVA6Cfg[579-:32]) >= 1 ? $clog2(CVA6Cfg[579-:32]) : 2 - $clog2(CVA6Cfg[579-:32]))) - 1)-:($clog2(CVA6Cfg[579-:32]) >= 1 ? $clog2(CVA6Cfg[579-:32]) : 2 - $clog2(CVA6Cfg[579-:32]))] * 2+:2]);
			// Trace: core/frontend/frontend.sv:181:5
			assign btb_prediction_shifted[0+:1 + CVA6Cfg[17070-:32]] = (serving_unaligned ? btb_q : btb_prediction[addr[0 + ($clog2(CVA6Cfg[579-:32]) >= 1 ? $clog2(CVA6Cfg[579-:32]) : ($clog2(CVA6Cfg[579-:32]) + ($clog2(CVA6Cfg[579-:32]) >= 1 ? $clog2(CVA6Cfg[579-:32]) : 2 - $clog2(CVA6Cfg[579-:32]))) - 1)-:($clog2(CVA6Cfg[579-:32]) >= 1 ? $clog2(CVA6Cfg[579-:32]) : 2 - $clog2(CVA6Cfg[579-:32]))] * (1 + CVA6Cfg[17070-:32])+:1 + CVA6Cfg[17070-:32]]);
			genvar _gv_i_17;
			for (_gv_i_17 = 1; _gv_i_17 < CVA6Cfg[579-:32]; _gv_i_17 = _gv_i_17 + 1) begin : gen_prediction_address
				localparam i = _gv_i_17;
				// Trace: core/frontend/frontend.sv:188:7
				assign bht_prediction_shifted[i * 2+:2] = bht_prediction[addr[(i * CVA6Cfg[17070-:32]) + ($clog2(CVA6Cfg[579-:32]) >= 1 ? $clog2(CVA6Cfg[579-:32]) : ($clog2(CVA6Cfg[579-:32]) + ($clog2(CVA6Cfg[579-:32]) >= 1 ? $clog2(CVA6Cfg[579-:32]) : 2 - $clog2(CVA6Cfg[579-:32]))) - 1)-:($clog2(CVA6Cfg[579-:32]) >= 1 ? $clog2(CVA6Cfg[579-:32]) : 2 - $clog2(CVA6Cfg[579-:32]))] * 2+:2];
				// Trace: core/frontend/frontend.sv:189:7
				assign btb_prediction_shifted[i * (1 + CVA6Cfg[17070-:32])+:1 + CVA6Cfg[17070-:32]] = btb_prediction[addr[(i * CVA6Cfg[17070-:32]) + ($clog2(CVA6Cfg[579-:32]) >= 1 ? $clog2(CVA6Cfg[579-:32]) : ($clog2(CVA6Cfg[579-:32]) + ($clog2(CVA6Cfg[579-:32]) >= 1 ? $clog2(CVA6Cfg[579-:32]) : 2 - $clog2(CVA6Cfg[579-:32]))) - 1)-:($clog2(CVA6Cfg[579-:32]) >= 1 ? $clog2(CVA6Cfg[579-:32]) : 2 - $clog2(CVA6Cfg[579-:32]))] * (1 + CVA6Cfg[17070-:32])+:1 + CVA6Cfg[17070-:32]];
			end
		end
		else begin : genblk2
			// Trace: core/frontend/frontend.sv:192:5
			assign bht_prediction_shifted[0+:2] = (serving_unaligned ? bht_q : bht_prediction[addr[1] * 2+:2]);
			// Trace: core/frontend/frontend.sv:193:5
			assign btb_prediction_shifted[0+:1 + CVA6Cfg[17070-:32]] = (serving_unaligned ? btb_q : btb_prediction[addr[1] * (1 + CVA6Cfg[17070-:32])+:1 + CVA6Cfg[17070-:32]]);
		end
	endgenerate
	// Trace: core/frontend/frontend.sv:199:3
	reg bp_valid;
	// Trace: core/frontend/frontend.sv:201:3
	wire [CVA6Cfg[579-:32] - 1:0] is_branch;
	// Trace: core/frontend/frontend.sv:202:3
	wire [CVA6Cfg[579-:32] - 1:0] is_call;
	// Trace: core/frontend/frontend.sv:203:3
	wire [CVA6Cfg[579-:32] - 1:0] is_jump;
	// Trace: core/frontend/frontend.sv:204:3
	wire [CVA6Cfg[579-:32] - 1:0] is_return;
	// Trace: core/frontend/frontend.sv:205:3
	wire [CVA6Cfg[579-:32] - 1:0] is_jalr;
	// Trace: core/frontend/frontend.sv:207:3
	genvar _gv_i_18;
	generate
		for (_gv_i_18 = 0; _gv_i_18 < CVA6Cfg[579-:32]; _gv_i_18 = _gv_i_18 + 1) begin : genblk3
			localparam i = _gv_i_18;
			// Trace: core/frontend/frontend.sv:209:5
			assign is_branch[i] = instruction_valid[i] & (rvi_branch[i] | rvc_branch[i]);
			// Trace: core/frontend/frontend.sv:211:5
			assign is_call[i] = instruction_valid[i] & (rvi_call[i] | rvc_call[i]);
			// Trace: core/frontend/frontend.sv:213:5
			assign is_return[i] = instruction_valid[i] & (rvi_return[i] | rvc_return[i]);
			// Trace: core/frontend/frontend.sv:215:5
			assign is_jump[i] = instruction_valid[i] & (rvi_jump[i] | rvc_jump[i]);
			// Trace: core/frontend/frontend.sv:217:5
			assign is_jalr[i] = (instruction_valid[i] & ~is_return[i]) & ((rvi_jalr[i] | rvc_jalr[i]) | rvc_jr[i]);
		end
	endgenerate
	// Trace: core/frontend/frontend.sv:221:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: core/frontend/frontend.sv:222:5
		taken_rvi_cf = 1'sb0;
		// Trace: core/frontend/frontend.sv:223:5
		taken_rvc_cf = 1'sb0;
		// Trace: core/frontend/frontend.sv:224:5
		predict_address = 1'sb0;
		// Trace: core/frontend/frontend.sv:226:5
		begin : sv2v_autoblock_1
			// Trace: core/frontend/frontend.sv:226:10
			reg signed [31:0] i;
			// Trace: core/frontend/frontend.sv:226:10
			for (i = 0; i < CVA6Cfg[579-:32]; i = i + 1)
				begin
					// Trace: core/frontend/frontend.sv:226:55
					cf_type[i * 3+:3] = 3'd0;
				end
		end
		// Trace: core/frontend/frontend.sv:228:5
		ras_push = 1'b0;
		// Trace: core/frontend/frontend.sv:229:5
		ras_pop = 1'b0;
		// Trace: core/frontend/frontend.sv:230:5
		ras_update = 1'sb0;
		begin : sv2v_autoblock_2
			// Trace: core/frontend/frontend.sv:233:10
			reg signed [31:0] i;
			// Trace: core/frontend/frontend.sv:233:10
			for (i = CVA6Cfg[579-:32] - 1; i >= 0; i = i - 1)
				begin
					// Trace: core/frontend/frontend.sv:234:7
					(* full_case, parallel_case *)
					case ({is_branch[i], is_return[i], is_jump[i], is_jalr[i]})
						4'b0000:
							;
						4'b0001: begin
							// Trace: core/frontend/frontend.sv:240:11
							ras_pop = 1'b0;
							// Trace: core/frontend/frontend.sv:241:11
							ras_push = 1'b0;
							// Trace: core/frontend/frontend.sv:242:11
							if (CVA6Cfg[16204-:32] && btb_prediction_shifted[(i * (1 + CVA6Cfg[17070-:32])) + (CVA6Cfg[17070-:32] + 0)]) begin
								// Trace: core/frontend/frontend.sv:243:13
								predict_address = btb_prediction_shifted[(i * (1 + CVA6Cfg[17070-:32])) + (CVA6Cfg[17070-:32] - 1)-:CVA6Cfg[17070-:32]];
								// Trace: core/frontend/frontend.sv:244:13
								cf_type[i * 3+:3] = 3'd3;
							end
						end
						4'b0010: begin
							// Trace: core/frontend/frontend.sv:249:11
							ras_pop = 1'b0;
							// Trace: core/frontend/frontend.sv:250:11
							ras_push = 1'b0;
							// Trace: core/frontend/frontend.sv:251:11
							taken_rvi_cf[i] = rvi_jump[i];
							// Trace: core/frontend/frontend.sv:252:11
							taken_rvc_cf[i] = rvc_jump[i];
							// Trace: core/frontend/frontend.sv:253:11
							cf_type[i * 3+:3] = 3'd2;
						end
						4'b0100: begin
							// Trace: core/frontend/frontend.sv:258:11
							ras_pop = ras_predict[CVA6Cfg[17070-:32] + 0] & instr_queue_consumed[i];
							// Trace: core/frontend/frontend.sv:259:11
							ras_push = 1'b0;
							// Trace: core/frontend/frontend.sv:260:11
							predict_address = ras_predict[CVA6Cfg[17070-:32] - 1-:CVA6Cfg[17070-:32]];
							// Trace: core/frontend/frontend.sv:261:11
							cf_type[i * 3+:3] = 3'd4;
						end
						4'b1000: begin
							// Trace: core/frontend/frontend.sv:265:11
							ras_pop = 1'b0;
							// Trace: core/frontend/frontend.sv:266:11
							ras_push = 1'b0;
							// Trace: core/frontend/frontend.sv:268:11
							if (bht_prediction_shifted[(i * 2) + 1]) begin
								// Trace: core/frontend/frontend.sv:269:13
								taken_rvi_cf[i] = rvi_branch[i] & bht_prediction_shifted[i * 2];
								// Trace: core/frontend/frontend.sv:270:13
								taken_rvc_cf[i] = rvc_branch[i] & bht_prediction_shifted[i * 2];
							end
							else begin
								// Trace: core/frontend/frontend.sv:274:13
								taken_rvi_cf[i] = rvi_branch[i] & rvi_imm[(i * CVA6Cfg[17070-:32]) + (CVA6Cfg[17070-:32] - 1)];
								// Trace: core/frontend/frontend.sv:275:13
								taken_rvc_cf[i] = rvc_branch[i] & rvc_imm[(i * CVA6Cfg[17070-:32]) + (CVA6Cfg[17070-:32] - 1)];
							end
							if (taken_rvi_cf[i] || taken_rvc_cf[i])
								// Trace: core/frontend/frontend.sv:278:13
								cf_type[i * 3+:3] = 3'd1;
						end
						default:
							;
					endcase
					if (is_call[i]) begin
						// Trace: core/frontend/frontend.sv:287:9
						ras_push = instr_queue_consumed[i];
						// Trace: core/frontend/frontend.sv:288:9
						ras_update = addr[i * CVA6Cfg[17070-:32]+:CVA6Cfg[17070-:32]] + (rvc_call[i] ? 2 : 4);
					end
					if (taken_rvc_cf[i] || taken_rvi_cf[i])
						// Trace: core/frontend/frontend.sv:292:9
						predict_address = addr[i * CVA6Cfg[17070-:32]+:CVA6Cfg[17070-:32]] + (taken_rvc_cf[i] ? rvc_imm[i * CVA6Cfg[17070-:32]+:CVA6Cfg[17070-:32]] : rvi_imm[i * CVA6Cfg[17070-:32]+:CVA6Cfg[17070-:32]]);
				end
		end
	end
	// Trace: core/frontend/frontend.sv:297:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: core/frontend/frontend.sv:298:5
		bp_valid = 1'b0;
		// Trace: core/frontend/frontend.sv:302:5
		begin : sv2v_autoblock_3
			// Trace: core/frontend/frontend.sv:302:10
			reg signed [31:0] i;
			// Trace: core/frontend/frontend.sv:302:10
			for (i = 0; i < CVA6Cfg[579-:32]; i = i + 1)
				begin
					// Trace: core/frontend/frontend.sv:303:5
					bp_valid = bp_valid | (((cf_type[i * 3+:3] != 3'd0) & (cf_type[i * 3+:3] != 3'd4)) | ((cf_type[i * 3+:3] == 3'd4) & ras_predict[CVA6Cfg[17070-:32] + 0]));
				end
		end
	end
	// Trace: core/frontend/frontend.sv:305:3
	assign is_mispredict = resolved_branch_i[1 + (bp_resolve_t_CVA6Cfg[9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (bp_resolve_t_CVA6Cfg[9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 4))] & resolved_branch_i[4];
	// Trace: core/frontend/frontend.sv:308:3
	wire [1:1] sv2v_tmp_32AF3;
	assign sv2v_tmp_32AF3 = instr_queue_ready;
	always @(*) icache_dreq_o[2 + (icache_dreq_t_CVA6Cfg[9509 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 1)] = sv2v_tmp_32AF3;
	// Trace: core/frontend/frontend.sv:309:3
	assign if_ready = icache_dreq_i[2 + (icache_drsp_t_CVA6Cfg[643-:32] + (icache_drsp_t_CVA6Cfg[708-:32] + (icache_drsp_t_CVA6Cfg[9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (((((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33) >= 0 ? ((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 34 : 1 - (((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33)) - 1))))] & instr_queue_ready;
	// Trace: core/frontend/frontend.sv:314:3
	wire [1:1] sv2v_tmp_C5596;
	assign sv2v_tmp_C5596 = (is_mispredict | flush_i) | replay;
	always @(*) icache_dreq_o[2 + (icache_dreq_t_CVA6Cfg[9509 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0)] = sv2v_tmp_C5596;
	// Trace: core/frontend/frontend.sv:317:3
	wire [1:1] sv2v_tmp_9A12C;
	assign sv2v_tmp_9A12C = icache_dreq_o[2 + (icache_dreq_t_CVA6Cfg[9509 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0)] | bp_valid;
	always @(*) icache_dreq_o[icache_dreq_t_CVA6Cfg[9509 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 1] = sv2v_tmp_9A12C;
	// Trace: core/frontend/frontend.sv:320:3
	wire [(1 + CVA6Cfg[17070-:32]) + 0:0] bht_update;
	// Trace: core/frontend/frontend.sv:321:3
	wire [((1 + CVA6Cfg[17070-:32]) + CVA6Cfg[17070-:32]) - 1:0] btb_update;
	// Trace: core/frontend/frontend.sv:324:3
	reg speculative_q;
	wire speculative_d;
	// Trace: core/frontend/frontend.sv:325:3
	assign speculative_d = ((((speculative_q && !resolved_branch_i[1 + (bp_resolve_t_CVA6Cfg[9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (bp_resolve_t_CVA6Cfg[9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 4))]) || |is_branch) || |is_return) || |is_jalr) && !flush_i;
	// Trace: core/frontend/frontend.sv:326:3
	wire [1:1] sv2v_tmp_9C044;
	assign sv2v_tmp_9C044 = speculative_d;
	always @(*) icache_dreq_o[icache_dreq_t_CVA6Cfg[9509 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0] = sv2v_tmp_9C044;
	// Trace: core/frontend/frontend.sv:328:3
	assign bht_update[1 + (CVA6Cfg[17070-:32] + 0)] = resolved_branch_i[1 + (bp_resolve_t_CVA6Cfg[9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (bp_resolve_t_CVA6Cfg[9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 4))] & (resolved_branch_i[2-:3] == 3'd1);
	// Trace: core/frontend/frontend.sv:330:3
	assign bht_update[CVA6Cfg[17070-:32] + 0-:((CVA6Cfg[17070-:32] + 0) >= 1 ? CVA6Cfg[17070-:32] + 0 : 2 - (CVA6Cfg[17070-:32] + 0))] = resolved_branch_i[bp_resolve_t_CVA6Cfg[9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (bp_resolve_t_CVA6Cfg[9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 4)-:((bp_resolve_t_CVA6Cfg[9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (bp_resolve_t_CVA6Cfg[9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 4)) >= (bp_resolve_t_CVA6Cfg[9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 5) ? ((bp_resolve_t_CVA6Cfg[9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (bp_resolve_t_CVA6Cfg[9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 4)) - (bp_resolve_t_CVA6Cfg[9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 5)) + 1 : ((bp_resolve_t_CVA6Cfg[9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 5) - (bp_resolve_t_CVA6Cfg[9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (bp_resolve_t_CVA6Cfg[9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 4))) + 1)];
	// Trace: core/frontend/frontend.sv:331:3
	assign bht_update[0] = resolved_branch_i[3];
	// Trace: core/frontend/frontend.sv:333:3
	assign btb_update[1 + (CVA6Cfg[17070-:32] + (CVA6Cfg[17070-:32] - 1))] = (resolved_branch_i[1 + (bp_resolve_t_CVA6Cfg[9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (bp_resolve_t_CVA6Cfg[9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 4))] & resolved_branch_i[4]) & (resolved_branch_i[2-:3] == 3'd3);
	// Trace: core/frontend/frontend.sv:336:3
	assign btb_update[CVA6Cfg[17070-:32] + (CVA6Cfg[17070-:32] - 1)-:((CVA6Cfg[17070-:32] + (CVA6Cfg[17070-:32] - 1)) >= (CVA6Cfg[17070-:32] + 0) ? ((CVA6Cfg[17070-:32] + (CVA6Cfg[17070-:32] - 1)) - (CVA6Cfg[17070-:32] + 0)) + 1 : ((CVA6Cfg[17070-:32] + 0) - (CVA6Cfg[17070-:32] + (CVA6Cfg[17070-:32] - 1))) + 1)] = resolved_branch_i[bp_resolve_t_CVA6Cfg[9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (bp_resolve_t_CVA6Cfg[9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 4)-:((bp_resolve_t_CVA6Cfg[9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (bp_resolve_t_CVA6Cfg[9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 4)) >= (bp_resolve_t_CVA6Cfg[9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 5) ? ((bp_resolve_t_CVA6Cfg[9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (bp_resolve_t_CVA6Cfg[9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 4)) - (bp_resolve_t_CVA6Cfg[9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 5)) + 1 : ((bp_resolve_t_CVA6Cfg[9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 5) - (bp_resolve_t_CVA6Cfg[9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (bp_resolve_t_CVA6Cfg[9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 4))) + 1)];
	// Trace: core/frontend/frontend.sv:337:3
	assign btb_update[CVA6Cfg[17070-:32] - 1-:CVA6Cfg[17070-:32]] = resolved_branch_i[bp_resolve_t_CVA6Cfg[9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 4-:((bp_resolve_t_CVA6Cfg[9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 4) >= 5 ? bp_resolve_t_CVA6Cfg[9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0 : 6 - (bp_resolve_t_CVA6Cfg[9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 4))];
	// Trace: core/frontend/frontend.sv:351:3
	always @(*) begin : npc_select
		// Trace: core/frontend/frontend.sv:352:5
		reg [CVA6Cfg[17070-:32] - 1:0] fetch_address;
		if (_sv2v_0)
			;
		// Trace: core/frontend/frontend.sv:359:5
		if (npc_rst_load_q) begin
			// Trace: core/frontend/frontend.sv:360:7
			npc_d = boot_addr_i;
			// Trace: core/frontend/frontend.sv:361:7
			fetch_address = boot_addr_i;
		end
		else begin
			// Trace: core/frontend/frontend.sv:363:7
			fetch_address = npc_q;
			// Trace: core/frontend/frontend.sv:365:7
			npc_d = npc_q;
		end
		if (bp_valid) begin
			// Trace: core/frontend/frontend.sv:369:7
			fetch_address = predict_address;
			// Trace: core/frontend/frontend.sv:370:7
			npc_d = predict_address;
		end
		if (if_ready)
			// Trace: core/frontend/frontend.sv:374:7
			npc_d = {fetch_address[CVA6Cfg[17070-:32] - 1:CVA6Cfg[611-:32]] + 1, {CVA6Cfg[611-:32] {1'b0}}};
		if (replay)
			// Trace: core/frontend/frontend.sv:380:7
			npc_d = replay_addr;
		if (is_mispredict)
			// Trace: core/frontend/frontend.sv:384:7
			npc_d = resolved_branch_i[bp_resolve_t_CVA6Cfg[9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 4-:((bp_resolve_t_CVA6Cfg[9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 4) >= 5 ? bp_resolve_t_CVA6Cfg[9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0 : 6 - (bp_resolve_t_CVA6Cfg[9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + (32 + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + ((bp_resolve_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 4))];
		if (eret_i)
			// Trace: core/frontend/frontend.sv:388:7
			npc_d = epc_i;
		if (ex_valid_i)
			// Trace: core/frontend/frontend.sv:392:7
			npc_d = trap_vector_base_i;
		if (set_pc_commit_i)
			// Trace: core/frontend/frontend.sv:404:7
			npc_d = pc_commit_i + (halt_i ? {CVA6Cfg[17070-:32] {1'sb0}} : {{CVA6Cfg[17070-:32] - 3 {1'b0}}, 3'b100});
		if (CVA6Cfg[1321] && set_debug_pc_i)
			// Trace: core/frontend/frontend.sv:409:7
			npc_d = CVA6Cfg[15915 + CVA6Cfg[17070-:32]:15916] + CVA6Cfg[16300 + CVA6Cfg[17070-:32]:16301];
		// Trace: core/frontend/frontend.sv:410:5
		icache_dreq_o[icache_dreq_t_CVA6Cfg[9509 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1-:icache_dreq_t_CVA6Cfg[9509 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + ((icache_dreq_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]] = fetch_address;
	end
	// Trace: core/frontend/frontend.sv:413:3
	wire [CVA6Cfg[643-:32] - 1:0] icache_data;
	// Trace: core/frontend/frontend.sv:415:3
	assign icache_data = icache_dreq_i[icache_drsp_t_CVA6Cfg[643-:32] + (icache_drsp_t_CVA6Cfg[708-:32] + (icache_drsp_t_CVA6Cfg[9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (((((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33) >= 0 ? ((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 34 : 1 - (((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33)) - 1)))-:((icache_drsp_t_CVA6Cfg[643-:32] + (icache_drsp_t_CVA6Cfg[708-:32] + (icache_drsp_t_CVA6Cfg[9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (((((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33) >= 0 ? ((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 34 : 1 - (((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33)) - 1)))) >= (icache_drsp_t_CVA6Cfg[708-:32] + (icache_drsp_t_CVA6Cfg[9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (((((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33) >= 0 ? ((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 34 : 1 - (((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33)) + 0))) ? ((icache_drsp_t_CVA6Cfg[643-:32] + (icache_drsp_t_CVA6Cfg[708-:32] + (icache_drsp_t_CVA6Cfg[9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (((((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33) >= 0 ? ((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 34 : 1 - (((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33)) - 1)))) - (icache_drsp_t_CVA6Cfg[708-:32] + (icache_drsp_t_CVA6Cfg[9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (((((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33) >= 0 ? ((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 34 : 1 - (((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33)) + 0)))) + 1 : ((icache_drsp_t_CVA6Cfg[708-:32] + (icache_drsp_t_CVA6Cfg[9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (((((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33) >= 0 ? ((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 34 : 1 - (((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33)) + 0))) - (icache_drsp_t_CVA6Cfg[643-:32] + (icache_drsp_t_CVA6Cfg[708-:32] + (icache_drsp_t_CVA6Cfg[9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (((((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33) >= 0 ? ((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 34 : 1 - (((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33)) - 1))))) + 1)] >> {shamt, 4'b0000};
	// Trace: core/frontend/frontend.sv:417:3
	localparam cva6_config_pkg_CVA6ConfigXlen = 64;
	localparam riscv_XLEN = cva6_config_pkg_CVA6ConfigXlen;
	localparam [63:0] riscv_INSTR_ACCESS_FAULT = 1;
	localparam [63:0] riscv_INSTR_GUEST_PAGE_FAULT = 20;
	localparam [63:0] riscv_INSTR_PAGE_FAULT = 12;
	always @(posedge clk_i or negedge rst_ni)
		// Trace: core/frontend/frontend.sv:418:5
		if (!rst_ni) begin
			// Trace: core/frontend/frontend.sv:419:7
			npc_rst_load_q <= 1'b1;
			// Trace: core/frontend/frontend.sv:420:7
			npc_q <= 1'sb0;
			// Trace: core/frontend/frontend.sv:421:7
			speculative_q <= 1'sb0;
			// Trace: core/frontend/frontend.sv:422:7
			icache_data_q <= 1'sb0;
			// Trace: core/frontend/frontend.sv:423:7
			icache_valid_q <= 1'b0;
			// Trace: core/frontend/frontend.sv:424:7
			icache_vaddr_q <= 'b0;
			// Trace: core/frontend/frontend.sv:425:7
			icache_gpaddr_q <= 'b0;
			// Trace: core/frontend/frontend.sv:426:7
			icache_tinst_q <= 'b0;
			// Trace: core/frontend/frontend.sv:427:7
			icache_gva_q <= 1'b0;
			// Trace: core/frontend/frontend.sv:428:7
			icache_ex_valid_q <= 2'd0;
			// Trace: core/frontend/frontend.sv:429:7
			btb_q <= 1'sb0;
			// Trace: core/frontend/frontend.sv:430:7
			bht_q <= 1'sb0;
		end
		else begin
			// Trace: core/frontend/frontend.sv:432:7
			npc_rst_load_q <= 1'b0;
			// Trace: core/frontend/frontend.sv:433:7
			npc_q <= npc_d;
			// Trace: core/frontend/frontend.sv:434:7
			speculative_q <= speculative_d;
			// Trace: core/frontend/frontend.sv:435:7
			icache_valid_q <= icache_dreq_i[1 + (icache_drsp_t_CVA6Cfg[643-:32] + (icache_drsp_t_CVA6Cfg[708-:32] + (icache_drsp_t_CVA6Cfg[9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (((((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33) >= 0 ? ((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 34 : 1 - (((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33)) - 1))))];
			// Trace: core/frontend/frontend.sv:436:7
			if (icache_dreq_i[1 + (icache_drsp_t_CVA6Cfg[643-:32] + (icache_drsp_t_CVA6Cfg[708-:32] + (icache_drsp_t_CVA6Cfg[9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (((((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33) >= 0 ? ((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 34 : 1 - (((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33)) - 1))))]) begin
				// Trace: core/frontend/frontend.sv:437:9
				icache_data_q <= icache_data;
				// Trace: core/frontend/frontend.sv:438:9
				icache_vaddr_q <= icache_dreq_i[icache_drsp_t_CVA6Cfg[9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (((((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33) >= 0 ? ((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 34 : 1 - (((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33)) - 1)-:((icache_drsp_t_CVA6Cfg[9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (((((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33) >= 0 ? ((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 34 : 1 - (((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33)) - 1)) >= (((((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33) >= 0 ? ((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 34 : 1 - (((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33)) + 0) ? ((icache_drsp_t_CVA6Cfg[9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (((((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33) >= 0 ? ((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 34 : 1 - (((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33)) - 1)) - (((((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33) >= 0 ? ((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 34 : 1 - (((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33)) + 0)) + 1 : ((((((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33) >= 0 ? ((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 34 : 1 - (((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33)) + 0) - (icache_drsp_t_CVA6Cfg[9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (((((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33) >= 0 ? ((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 34 : 1 - (((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33)) - 1))) + 1)];
				// Trace: core/frontend/frontend.sv:439:9
				if (CVA6Cfg[16543]) begin
					// Trace: core/frontend/frontend.sv:440:11
					icache_gpaddr_q <= icache_dreq_i[((((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33) >= 0 ? (((((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33) >= 0 ? ((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 34 : 1 - (((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33)) - 1) - ((((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33) - ((icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 33) - ((icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1) - (CVA6Cfg[17006-:32] - 1)))) : 0 + (((icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1) - (CVA6Cfg[17006-:32] - 1)) - (icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 33))):((((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33) >= 0 ? (((((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33) >= 0 ? ((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 34 : 1 - (((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33)) - 1) - ((((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33) - ((icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 33) - (icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1))) : 0 + ((icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1) - (icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 33)))];
					// Trace: core/frontend/frontend.sv:441:11
					icache_tinst_q <= icache_dreq_i[((((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33) >= 0 ? (((((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33) >= 0 ? ((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 34 : 1 - (((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33)) - 1) - (((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 0) : -2)-:32];
					// Trace: core/frontend/frontend.sv:442:11
					icache_gva_q <= icache_dreq_i[((((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33) >= 0 ? (((((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33) >= 0 ? ((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 34 : 1 - (((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33)) - 1) - (((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 32) : -1)];
				end
				else begin
					// Trace: core/frontend/frontend.sv:444:11
					icache_gpaddr_q <= 'b0;
					// Trace: core/frontend/frontend.sv:445:11
					icache_tinst_q <= 'b0;
					// Trace: core/frontend/frontend.sv:446:11
					icache_gva_q <= 1'b0;
				end
				if (CVA6Cfg[16367] && (icache_dreq_i[((((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33) >= 0 ? (((((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33) >= 0 ? ((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 34 : 1 - (((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33)) - 1) - ((((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33) - (icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 33)))) : (((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 33))) >= (icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 34)) ? ((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 33))) - (icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 34))) + 1 : ((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 34)) - (icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 33)))) + 1) - (icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 33)))) - 1)-:((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 33))) >= (icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 34)) ? ((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 33))) - (icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 34))) + 1 : ((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 34)) - (icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 33)))) + 1)] == riscv_INSTR_GUEST_PAGE_FAULT))
					// Trace: core/frontend/frontend.sv:451:11
					icache_ex_valid_q <= 2'd3;
				else if (CVA6Cfg[16367] && (icache_dreq_i[((((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33) >= 0 ? (((((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33) >= 0 ? ((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 34 : 1 - (((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33)) - 1) - ((((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33) - (icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 33)))) : (((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 33))) >= (icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 34)) ? ((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 33))) - (icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 34))) + 1 : ((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 34)) - (icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 33)))) + 1) - (icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 33)))) - 1)-:((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 33))) >= (icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 34)) ? ((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 33))) - (icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 34))) + 1 : ((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 34)) - (icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 33)))) + 1)] == riscv_INSTR_PAGE_FAULT))
					// Trace: core/frontend/frontend.sv:453:11
					icache_ex_valid_q <= 2'd2;
				else if (icache_dreq_i[((((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33) >= 0 ? (((((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33) >= 0 ? ((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 34 : 1 - (((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33)) - 1) - ((((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33) - (icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 33)))) : (((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 33))) >= (icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 34)) ? ((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 33))) - (icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 34))) + 1 : ((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 34)) - (icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 33)))) + 1) - (icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 33)))) - 1)-:((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 33))) >= (icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 34)) ? ((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 33))) - (icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 34))) + 1 : ((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 34)) - (icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 33)))) + 1)] == riscv_INSTR_ACCESS_FAULT)
					// Trace: core/frontend/frontend.sv:455:11
					icache_ex_valid_q <= 2'd1;
				else
					// Trace: core/frontend/frontend.sv:457:11
					icache_ex_valid_q <= 2'd0;
				// Trace: core/frontend/frontend.sv:460:9
				btb_q <= btb_prediction[(CVA6Cfg[579-:32] - 1) * (1 + CVA6Cfg[17070-:32])+:1 + CVA6Cfg[17070-:32]];
				// Trace: core/frontend/frontend.sv:461:9
				bht_q <= bht_prediction[(CVA6Cfg[579-:32] - 1) * 2+:2];
			end
		end
	// Trace: core/frontend/frontend.sv:466:3
	generate
		if (CVA6Cfg[16236-:32] == 0) begin : genblk4
			// Trace: core/frontend/frontend.sv:467:5
			assign ras_predict = 1'sb0;
		end
		else begin : ras_gen
			// Trace: core/frontend/frontend.sv:469:5
			ras_091E3_171B5 #(
				.ras_t_CVA6Cfg(CVA6Cfg),
				.ras_t_config_pkg_NrMaxRules(config_pkg_NrMaxRules),
				.CVA6Cfg(CVA6Cfg),
				.DEPTH(CVA6Cfg[16236-:32])
			) i_ras(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.flush_bp_i(flush_bp_i),
				.push_i(ras_push),
				.pop_i(ras_pop),
				.data_i(ras_update),
				.data_o(ras_predict)
			);
		end
	endgenerate
	// Trace: core/frontend/frontend.sv:487:3
	assign vpc_btb = (CVA6Cfg[16876] ? icache_dreq_i[icache_drsp_t_CVA6Cfg[9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (((((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33) >= 0 ? ((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 34 : 1 - (((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33)) - 1)-:((icache_drsp_t_CVA6Cfg[9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (((((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33) >= 0 ? ((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 34 : 1 - (((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33)) - 1)) >= (((((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33) >= 0 ? ((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 34 : 1 - (((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33)) + 0) ? ((icache_drsp_t_CVA6Cfg[9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (((((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33) >= 0 ? ((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 34 : 1 - (((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33)) - 1)) - (((((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33) >= 0 ? ((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 34 : 1 - (((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33)) + 0)) + 1 : ((((((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33) >= 0 ? ((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 34 : 1 - (((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33)) + 0) - (icache_drsp_t_CVA6Cfg[9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (((((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33) >= 0 ? ((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 34 : 1 - (((icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + icache_drsp_t_CVA6Cfg[9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + icache_drsp_t_CVA6Cfg[9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9413 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9445 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + (32 + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + ((icache_drsp_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 33)) - 1))) + 1)] : icache_vaddr_q);
	// Trace: core/frontend/frontend.sv:489:3
	generate
		if (CVA6Cfg[16204-:32] == 0) begin : genblk5
			// Trace: core/frontend/frontend.sv:490:5
			assign btb_prediction = 1'sb0;
		end
		else begin : btb_gen
			// Trace: core/frontend/frontend.sv:492:5
			btb_C3780_5CA66 #(
				.btb_prediction_t_CVA6Cfg(CVA6Cfg),
				.btb_prediction_t_config_pkg_NrMaxRules(config_pkg_NrMaxRules),
				.btb_update_t_CVA6Cfg(CVA6Cfg),
				.btb_update_t_config_pkg_NrMaxRules(config_pkg_NrMaxRules),
				.CVA6Cfg(CVA6Cfg),
				.NR_ENTRIES(CVA6Cfg[16204-:32])
			) i_btb(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.flush_bp_i(flush_bp_i),
				.debug_mode_i(debug_mode_i),
				.vpc_i(vpc_btb),
				.btb_update_i(btb_update),
				.btb_prediction_o(btb_prediction)
			);
		end
	endgenerate
	// Trace: core/frontend/frontend.sv:508:3
	generate
		if (CVA6Cfg[16172-:32] == 0) begin : genblk6
			// Trace: core/frontend/frontend.sv:509:5
			assign bht_prediction = 1'sb0;
		end
		else begin : bht_gen
			// Trace: core/frontend/frontend.sv:511:5
			bht_980B8_E74A8 #(
				.bht_update_t_CVA6Cfg(CVA6Cfg),
				.bht_update_t_config_pkg_NrMaxRules(config_pkg_NrMaxRules),
				.CVA6Cfg(CVA6Cfg),
				.NR_ENTRIES(CVA6Cfg[16172-:32])
			) i_bht(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.flush_bp_i(flush_bp_i),
				.debug_mode_i(debug_mode_i),
				.vpc_i(icache_vaddr_q),
				.bht_update_i(bht_update),
				.bht_prediction_o(bht_prediction)
			);
		end
	endgenerate
	// Trace: core/frontend/frontend.sv:528:3
	genvar _gv_i_19;
	generate
		for (_gv_i_19 = 0; _gv_i_19 < CVA6Cfg[579-:32]; _gv_i_19 = _gv_i_19 + 1) begin : gen_instr_scan
			localparam i = _gv_i_19;
			// Trace: core/frontend/frontend.sv:529:5
			instr_scan #(.CVA6Cfg(CVA6Cfg)) i_instr_scan(
				.instr_i(instr[i * 32+:32]),
				.rvi_return_o(rvi_return[i]),
				.rvi_call_o(rvi_call[i]),
				.rvi_branch_o(rvi_branch[i]),
				.rvi_jalr_o(rvi_jalr[i]),
				.rvi_jump_o(rvi_jump[i]),
				.rvi_imm_o(rvi_imm[i * CVA6Cfg[17070-:32]+:CVA6Cfg[17070-:32]]),
				.rvc_branch_o(rvc_branch[i]),
				.rvc_jump_o(rvc_jump[i]),
				.rvc_jr_o(rvc_jr[i]),
				.rvc_return_o(rvc_return[i]),
				.rvc_jalr_o(rvc_jalr[i]),
				.rvc_call_o(rvc_call[i]),
				.rvc_imm_o(rvc_imm[i * CVA6Cfg[17070-:32]+:CVA6Cfg[17070-:32]])
			);
		end
	endgenerate
	// Trace: core/frontend/frontend.sv:549:3
	instr_queue_F2351_A36A8 #(
		.fetch_entry_t_fetch_entry_t_CVA6Cfg(fetch_entry_t_CVA6Cfg),
		.fetch_entry_t_fetch_entry_t_config_pkg_NrMaxRules(fetch_entry_t_config_pkg_NrMaxRules),
		.CVA6Cfg(CVA6Cfg)
	) i_instr_queue(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(flush_i),
		.instr_i(instr),
		.addr_i(addr),
		.exception_i(icache_ex_valid_q),
		.exception_addr_i(icache_vaddr_q),
		.exception_gpaddr_i(icache_gpaddr_q),
		.exception_tinst_i(icache_tinst_q),
		.exception_gva_i(icache_gva_q),
		.predict_address_i(predict_address),
		.cf_type_i(cf_type),
		.valid_i(instruction_valid),
		.consumed_o(instr_queue_consumed),
		.ready_o(instr_queue_ready),
		.replay_o(replay),
		.replay_addr_o(replay_addr),
		.fetch_entry_o(fetch_entry_o),
		.fetch_entry_valid_o(fetch_entry_valid_o),
		.fetch_entry_ready_i(fetch_entry_ready_i)
	);
	// Trace: core/frontend/frontend.sv:577:3
	initial _sv2v_0 = 0;
endmodule
