// removed module with interface ports: axi_slice_wrap
