module fpnew_top_D81B0_8D9C0 (
	clk_i,
	rst_ni,
	operands_i,
	rnd_mode_i,
	op_i,
	op_mod_i,
	src_fmt_i,
	dst_fmt_i,
	int_fmt_i,
	vectorial_op_i,
	tag_i,
	simd_mask_i,
	in_valid_i,
	in_ready_o,
	flush_i,
	result_o,
	status_o,
	tag_o,
	out_valid_o,
	out_ready_i,
	busy_o
);
	// removed localparam type TagType_CVA6Cfg_type
	// removed localparam type TagType_config_pkg_NrMaxRules_type
	parameter [17102:0] TagType_CVA6Cfg = 0;
	parameter signed [31:0] TagType_config_pkg_NrMaxRules = 0;
	reg _sv2v_0;
	// Trace: core/cvfpu/src/fpnew_top.sv:18:13
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	// removed localparam type fpnew_pkg_fmt_logic_t
	localparam [31:0] fpnew_pkg_NUM_INT_FORMATS = 4;
	// removed localparam type fpnew_pkg_ifmt_logic_t
	// removed localparam type fpnew_pkg_fpu_features_t
	localparam [42:0] fpnew_pkg_RV64D_Xsflt = 43'h000000207ff;
	parameter [42:0] Features = fpnew_pkg_RV64D_Xsflt;
	// Trace: core/cvfpu/src/fpnew_top.sv:19:13
	// removed localparam type fpnew_pkg_pipe_config_t
	// removed localparam type fpnew_pkg_unit_type_t
	localparam [31:0] fpnew_pkg_NUM_OPGROUPS = 4;
	// removed localparam type fpnew_pkg_fmt_unit_types_t
	// removed localparam type fpnew_pkg_opgrp_fmt_unit_types_t
	// removed localparam type fpnew_pkg_fmt_unsigned_t
	// removed localparam type fpnew_pkg_opgrp_fmt_unsigned_t
	// removed localparam type fpnew_pkg_fpu_implementation_t
	function automatic [159:0] sv2v_cast_C3475;
		input reg [159:0] inp;
		sv2v_cast_C3475 = inp;
	endfunction
	function automatic [((32'd4 * 32'd5) * 32) - 1:0] sv2v_cast_52F10;
		input reg [((32'd4 * 32'd5) * 32) - 1:0] inp;
		sv2v_cast_52F10 = inp;
	endfunction
	function automatic [((32'd4 * 32'd5) * 2) - 1:0] sv2v_cast_18D94;
		input reg [((32'd4 * 32'd5) * 2) - 1:0] inp;
		sv2v_cast_18D94 = inp;
	endfunction
	localparam [(((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 32) + ((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 2)) + 1:0] fpnew_pkg_DEFAULT_NOREGS = {sv2v_cast_52F10({fpnew_pkg_NUM_OPGROUPS {sv2v_cast_C3475(0)}}), sv2v_cast_18D94({{fpnew_pkg_NUM_FP_FORMATS {2'd1}}, {fpnew_pkg_NUM_FP_FORMATS {2'd2}}, {fpnew_pkg_NUM_FP_FORMATS {2'd1}}, {fpnew_pkg_NUM_FP_FORMATS {2'd2}}}), 2'd0};
	parameter [(((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 32) + ((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 2)) + 1:0] Implementation = fpnew_pkg_DEFAULT_NOREGS;
	// Trace: core/cvfpu/src/fpnew_top.sv:20:45
	// removed localparam type TagType
	// Trace: core/cvfpu/src/fpnew_top.sv:21:13
	parameter [31:0] TrueSIMDClass = 0;
	// Trace: core/cvfpu/src/fpnew_top.sv:22:13
	parameter [31:0] EnableSIMDMask = 0;
	// Trace: core/cvfpu/src/fpnew_top.sv:24:14
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	// removed localparam type fpnew_pkg_fp_format_e
	// removed localparam type fpnew_pkg_fp_encoding_t
	localparam [319:0] fpnew_pkg_FP_ENCODINGS = 320'h8000000170000000b00000034000000050000000a00000005000000020000000800000007;
	function automatic [31:0] fpnew_pkg_fp_width;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:304:44
		input reg [2:0] fmt;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:305:5
		fpnew_pkg_fp_width = (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] + fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32]) + 1;
	endfunction
	function automatic signed [31:0] fpnew_pkg_maximum;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:296:34
		input reg signed [31:0] a;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:296:41
		input reg signed [31:0] b;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:297:5
		fpnew_pkg_maximum = (a > b ? a : b);
	endfunction
	function automatic [2:0] sv2v_cast_5D882;
		input reg [2:0] inp;
		sv2v_cast_5D882 = inp;
	endfunction
	function automatic [31:0] fpnew_pkg_max_fp_width;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:309:48
		input reg [0:4] cfg;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:310:5
		reg [31:0] res;
		begin
			res = 0;
			// Trace: core/cvfpu/src/fpnew_pkg.sv:311:5
			begin : sv2v_autoblock_1
				// Trace: core/cvfpu/src/fpnew_pkg.sv:311:10
				reg [31:0] i;
				// Trace: core/cvfpu/src/fpnew_pkg.sv:311:10
				for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
					if (cfg[i])
						// Trace: core/cvfpu/src/fpnew_pkg.sv:313:9
						res = $unsigned(fpnew_pkg_maximum(res, fpnew_pkg_fp_width(sv2v_cast_5D882(i))));
			end
			fpnew_pkg_max_fp_width = res;
		end
	endfunction
	function automatic signed [31:0] fpnew_pkg_minimum;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:292:34
		input reg signed [31:0] a;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:292:41
		input reg signed [31:0] b;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:293:5
		fpnew_pkg_minimum = (a < b ? a : b);
	endfunction
	function automatic [31:0] fpnew_pkg_min_fp_width;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:318:48
		input reg [0:4] cfg;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:319:5
		reg [31:0] res;
		begin
			res = fpnew_pkg_max_fp_width(cfg);
			// Trace: core/cvfpu/src/fpnew_pkg.sv:320:5
			begin : sv2v_autoblock_2
				// Trace: core/cvfpu/src/fpnew_pkg.sv:320:10
				reg [31:0] i;
				// Trace: core/cvfpu/src/fpnew_pkg.sv:320:10
				for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
					if (cfg[i])
						// Trace: core/cvfpu/src/fpnew_pkg.sv:322:9
						res = $unsigned(fpnew_pkg_minimum(res, fpnew_pkg_fp_width(sv2v_cast_5D882(i))));
			end
			fpnew_pkg_min_fp_width = res;
		end
	endfunction
	function automatic [31:0] fpnew_pkg_max_num_lanes;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:395:49
		input reg [31:0] width;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:395:69
		input reg [0:4] cfg;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:395:86
		input reg vec;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:396:5
		fpnew_pkg_max_num_lanes = (vec ? width / fpnew_pkg_min_fp_width(cfg) : 1);
	endfunction
	localparam [31:0] NumLanes = fpnew_pkg_max_num_lanes(Features[42-:32], Features[8-:5], Features[10]);
	// Trace: core/cvfpu/src/fpnew_top.sv:25:27
	// removed localparam type MaskType
	// Trace: core/cvfpu/src/fpnew_top.sv:26:14
	localparam [31:0] WIDTH = Features[42-:32];
	// Trace: core/cvfpu/src/fpnew_top.sv:27:14
	localparam [31:0] NUM_OPERANDS = 3;
	// Trace: core/cvfpu/src/fpnew_top.sv:29:3
	input wire clk_i;
	// Trace: core/cvfpu/src/fpnew_top.sv:30:3
	input wire rst_ni;
	// Trace: core/cvfpu/src/fpnew_top.sv:32:3
	input wire [(NUM_OPERANDS * WIDTH) - 1:0] operands_i;
	// Trace: core/cvfpu/src/fpnew_top.sv:33:3
	// removed localparam type fpnew_pkg_roundmode_e
	input wire [2:0] rnd_mode_i;
	// Trace: core/cvfpu/src/fpnew_top.sv:34:3
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	// removed localparam type fpnew_pkg_operation_e
	input wire [3:0] op_i;
	// Trace: core/cvfpu/src/fpnew_top.sv:35:3
	input wire op_mod_i;
	// Trace: core/cvfpu/src/fpnew_top.sv:36:3
	input wire [2:0] src_fmt_i;
	// Trace: core/cvfpu/src/fpnew_top.sv:37:3
	input wire [2:0] dst_fmt_i;
	// Trace: core/cvfpu/src/fpnew_top.sv:38:3
	localparam [31:0] fpnew_pkg_INT_FORMAT_BITS = 2;
	// removed localparam type fpnew_pkg_int_format_e
	input wire [1:0] int_fmt_i;
	// Trace: core/cvfpu/src/fpnew_top.sv:39:3
	input wire vectorial_op_i;
	// Trace: core/cvfpu/src/fpnew_top.sv:40:3
	input wire [TagType_CVA6Cfg[8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1:0] tag_i;
	// Trace: core/cvfpu/src/fpnew_top.sv:41:3
	input wire [NumLanes - 1:0] simd_mask_i;
	// Trace: core/cvfpu/src/fpnew_top.sv:43:3
	input wire in_valid_i;
	// Trace: core/cvfpu/src/fpnew_top.sv:44:3
	output wire in_ready_o;
	// Trace: core/cvfpu/src/fpnew_top.sv:45:3
	input wire flush_i;
	// Trace: core/cvfpu/src/fpnew_top.sv:47:3
	output wire [WIDTH - 1:0] result_o;
	// Trace: core/cvfpu/src/fpnew_top.sv:48:3
	// removed localparam type fpnew_pkg_status_t
	output wire [4:0] status_o;
	// Trace: core/cvfpu/src/fpnew_top.sv:49:3
	output wire [TagType_CVA6Cfg[8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1:0] tag_o;
	// Trace: core/cvfpu/src/fpnew_top.sv:51:3
	output wire out_valid_o;
	// Trace: core/cvfpu/src/fpnew_top.sv:52:3
	input wire out_ready_i;
	// Trace: core/cvfpu/src/fpnew_top.sv:54:3
	output wire busy_o;
	// Trace: core/cvfpu/src/fpnew_top.sv:57:3
	localparam [31:0] NUM_OPGROUPS = fpnew_pkg_NUM_OPGROUPS;
	// Trace: core/cvfpu/src/fpnew_top.sv:58:3
	localparam [31:0] NUM_FORMATS = fpnew_pkg_NUM_FP_FORMATS;
	// Trace: core/cvfpu/src/fpnew_top.sv:63:3
	// removed localparam type output_t
	// Trace: core/cvfpu/src/fpnew_top.sv:70:3
	wire [3:0] opgrp_in_ready;
	wire [3:0] opgrp_out_valid;
	wire [3:0] opgrp_out_ready;
	wire [3:0] opgrp_ext;
	wire [3:0] opgrp_busy;
	// Trace: core/cvfpu/src/fpnew_top.sv:71:3
	wire [(4 * ((WIDTH + 5) + TagType_CVA6Cfg[8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)])) - 1:0] opgrp_outputs;
	// Trace: core/cvfpu/src/fpnew_top.sv:73:3
	wire [(NUM_FORMATS * NUM_OPERANDS) - 1:0] is_boxed;
	// Trace: core/cvfpu/src/fpnew_top.sv:78:3
	// removed localparam type fpnew_pkg_opgroup_e
	function automatic [3:0] sv2v_cast_4CD2E;
		input reg [3:0] inp;
		sv2v_cast_4CD2E = inp;
	endfunction
	function automatic [1:0] fpnew_pkg_get_opgroup;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:368:44
		input reg [3:0] op;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:369:5
		(* full_case, parallel_case *)
		case (op)
			sv2v_cast_4CD2E(0), sv2v_cast_4CD2E(1), sv2v_cast_4CD2E(2), sv2v_cast_4CD2E(3): fpnew_pkg_get_opgroup = 2'd0;
			sv2v_cast_4CD2E(4), sv2v_cast_4CD2E(5): fpnew_pkg_get_opgroup = 2'd1;
			sv2v_cast_4CD2E(6), sv2v_cast_4CD2E(7), sv2v_cast_4CD2E(8), sv2v_cast_4CD2E(9): fpnew_pkg_get_opgroup = 2'd2;
			sv2v_cast_4CD2E(10), sv2v_cast_4CD2E(11), sv2v_cast_4CD2E(12), sv2v_cast_4CD2E(13), sv2v_cast_4CD2E(14): fpnew_pkg_get_opgroup = 2'd3;
			default: fpnew_pkg_get_opgroup = 2'd2;
		endcase
	endfunction
	assign in_ready_o = in_valid_i & opgrp_in_ready[fpnew_pkg_get_opgroup(op_i)];
	// Trace: core/cvfpu/src/fpnew_top.sv:81:3
	genvar _gv_fmt_12;
	function automatic signed [31:0] sv2v_cast_32_signed;
		input reg signed [31:0] inp;
		sv2v_cast_32_signed = inp;
	endfunction
	generate
		for (_gv_fmt_12 = 0; _gv_fmt_12 < sv2v_cast_32_signed(NUM_FORMATS); _gv_fmt_12 = _gv_fmt_12 + 1) begin : gen_nanbox_check
			localparam fmt = _gv_fmt_12;
			// Trace: core/cvfpu/src/fpnew_top.sv:82:5
			localparam [31:0] FP_WIDTH = fpnew_pkg_fp_width(sv2v_cast_5D882(fmt));
			if (Features[9] && (FP_WIDTH < WIDTH)) begin : check
				genvar _gv_op_3;
				for (_gv_op_3 = 0; _gv_op_3 < sv2v_cast_32_signed(NUM_OPERANDS); _gv_op_3 = _gv_op_3 + 1) begin : operands
					localparam op = _gv_op_3;
					// Trace: core/cvfpu/src/fpnew_top.sv:86:9
					assign is_boxed[(fmt * NUM_OPERANDS) + op] = (!vectorial_op_i ? operands_i[(op * WIDTH) + ((WIDTH - 1) >= FP_WIDTH ? WIDTH - 1 : ((WIDTH - 1) + ((WIDTH - 1) >= FP_WIDTH ? ((WIDTH - 1) - FP_WIDTH) + 1 : (FP_WIDTH - (WIDTH - 1)) + 1)) - 1)-:((WIDTH - 1) >= FP_WIDTH ? ((WIDTH - 1) - FP_WIDTH) + 1 : (FP_WIDTH - (WIDTH - 1)) + 1)] == {((WIDTH - 1) >= FP_WIDTH ? ((WIDTH - 1) - FP_WIDTH) + 1 : (FP_WIDTH - (WIDTH - 1)) + 1) * 1 {1'sb1}} : 1'b1);
				end
			end
			else begin : no_check
				// Trace: core/cvfpu/src/fpnew_top.sv:91:7
				assign is_boxed[fmt * NUM_OPERANDS+:NUM_OPERANDS] = 1'sb1;
			end
		end
	endgenerate
	// Trace: core/cvfpu/src/fpnew_top.sv:96:3
	wire [NumLanes - 1:0] simd_mask;
	// Trace: core/cvfpu/src/fpnew_top.sv:97:3
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	assign simd_mask = simd_mask_i | ~{NumLanes {sv2v_cast_1(EnableSIMDMask)}};
	// Trace: core/cvfpu/src/fpnew_top.sv:102:3
	genvar _gv_opgrp_1;
	function automatic [31:0] fpnew_pkg_num_operands;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:379:48
		input reg [1:0] grp;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:380:5
		(* full_case, parallel_case *)
		case (grp)
			2'd0: fpnew_pkg_num_operands = 3;
			2'd1: fpnew_pkg_num_operands = 2;
			2'd2: fpnew_pkg_num_operands = 2;
			2'd3: fpnew_pkg_num_operands = 3;
			default: fpnew_pkg_num_operands = 0;
		endcase
	endfunction
	function automatic [1:0] sv2v_cast_2;
		input reg [1:0] inp;
		sv2v_cast_2 = inp;
	endfunction
	generate
		for (_gv_opgrp_1 = 0; _gv_opgrp_1 < sv2v_cast_32_signed(NUM_OPGROUPS); _gv_opgrp_1 = _gv_opgrp_1 + 1) begin : gen_operation_groups
			localparam opgrp = _gv_opgrp_1;
			// Trace: core/cvfpu/src/fpnew_top.sv:103:5
			localparam [31:0] NUM_OPS = fpnew_pkg_num_operands(sv2v_cast_2(opgrp));
			// Trace: core/cvfpu/src/fpnew_top.sv:105:5
			wire in_valid;
			// Trace: core/cvfpu/src/fpnew_top.sv:106:5
			reg [(NUM_FORMATS * NUM_OPS) - 1:0] input_boxed;
			// Trace: core/cvfpu/src/fpnew_top.sv:108:5
			assign in_valid = in_valid_i & (fpnew_pkg_get_opgroup(op_i) == sv2v_cast_2(opgrp));
			// Trace: core/cvfpu/src/fpnew_top.sv:111:5
			always @(*) begin : slice_inputs
				if (_sv2v_0)
					;
				// Trace: core/cvfpu/src/fpnew_top.sv:112:7
				begin : sv2v_autoblock_3
					// Trace: core/cvfpu/src/fpnew_top.sv:112:12
					reg [31:0] fmt;
					// Trace: core/cvfpu/src/fpnew_top.sv:112:12
					for (fmt = 0; fmt < NUM_FORMATS; fmt = fmt + 1)
						begin
							// Trace: core/cvfpu/src/fpnew_top.sv:113:9
							input_boxed[fmt * fpnew_pkg_num_operands(sv2v_cast_2(_gv_opgrp_1))+:fpnew_pkg_num_operands(sv2v_cast_2(_gv_opgrp_1))] = is_boxed[(fmt * NUM_OPERANDS) + (NUM_OPS - 1)-:NUM_OPS];
						end
				end
			end
			// Trace: core/cvfpu/src/fpnew_top.sv:116:5
			fpnew_opgroup_block_D3AB0_1C1E0 #(
				.TagType_TagType_CVA6Cfg(TagType_CVA6Cfg),
				.TagType_TagType_config_pkg_NrMaxRules(TagType_config_pkg_NrMaxRules),
				.OpGroup(sv2v_cast_2(opgrp)),
				.Width(WIDTH),
				.EnableVectors(Features[10]),
				.FpFmtMask(Features[8-:5]),
				.IntFmtMask(Features[3-:fpnew_pkg_NUM_INT_FORMATS]),
				.FmtPipeRegs(Implementation[(((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 32) + (((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 2) + 1)) - ((((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 32) - 1) - (32 * ((3 - opgrp) * fpnew_pkg_NUM_FP_FORMATS)))+:160]),
				.FmtUnitTypes(Implementation[(((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 2) + 1) - ((((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 2) - 1) - (2 * ((3 - opgrp) * fpnew_pkg_NUM_FP_FORMATS)))+:10]),
				.PipeConfig(Implementation[1-:2]),
				.TrueSIMDClass(TrueSIMDClass)
			) i_opgroup_block(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.operands_i(operands_i[WIDTH * ((NUM_OPS - 1) - (NUM_OPS - 1))+:WIDTH * NUM_OPS]),
				.is_boxed_i(input_boxed),
				.rnd_mode_i(rnd_mode_i),
				.op_i(op_i),
				.op_mod_i(op_mod_i),
				.src_fmt_i(src_fmt_i),
				.dst_fmt_i(dst_fmt_i),
				.int_fmt_i(int_fmt_i),
				.vectorial_op_i(vectorial_op_i),
				.tag_i(tag_i),
				.simd_mask_i(simd_mask),
				.in_valid_i(in_valid),
				.in_ready_o(opgrp_in_ready[opgrp]),
				.flush_i(flush_i),
				.result_o(opgrp_outputs[(opgrp * ((WIDTH + 5) + TagType_CVA6Cfg[8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)])) + (WIDTH + (TagType_CVA6Cfg[8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 4))-:((WIDTH + (TagType_CVA6Cfg[8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 4)) >= (5 + (TagType_CVA6Cfg[8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0)) ? ((WIDTH + (TagType_CVA6Cfg[8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 4)) - (5 + (TagType_CVA6Cfg[8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0))) + 1 : ((5 + (TagType_CVA6Cfg[8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0)) - (WIDTH + (TagType_CVA6Cfg[8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 4))) + 1)]),
				.status_o(opgrp_outputs[(opgrp * ((WIDTH + 5) + TagType_CVA6Cfg[8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)])) + (TagType_CVA6Cfg[8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 4)-:((TagType_CVA6Cfg[8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 4) >= (TagType_CVA6Cfg[8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0) ? ((TagType_CVA6Cfg[8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 4) - (TagType_CVA6Cfg[8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0)) + 1 : ((TagType_CVA6Cfg[8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0) - (TagType_CVA6Cfg[8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 4)) + 1)]),
				.extension_bit_o(opgrp_ext[opgrp]),
				.tag_o(opgrp_outputs[(opgrp * ((WIDTH + 5) + TagType_CVA6Cfg[8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)])) + (TagType_CVA6Cfg[8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1)-:TagType_CVA6Cfg[8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]]),
				.out_valid_o(opgrp_out_valid[opgrp]),
				.out_ready_i(opgrp_out_ready[opgrp]),
				.busy_o(opgrp_busy[opgrp])
			);
		end
	endgenerate
	// Trace: core/cvfpu/src/fpnew_top.sv:157:3
	wire [((WIDTH + 5) + TagType_CVA6Cfg[8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) - 1:0] arbiter_output;
	// Trace: core/cvfpu/src/fpnew_top.sv:160:3
	localparam [31:0] sv2v_uu_i_arbiter_NumIn = NUM_OPGROUPS;
	localparam [31:0] sv2v_uu_i_arbiter_IdxWidth = $unsigned(2);
	// removed localparam type sv2v_uu_i_arbiter_rr_i
	localparam [sv2v_uu_i_arbiter_IdxWidth - 1:0] sv2v_uu_i_arbiter_ext_rr_i_0 = 1'sb0;
	rr_arb_tree_1227C_AFDD0 #(
		.DataType_TagType_CVA6Cfg(TagType_CVA6Cfg),
		.DataType_TagType_config_pkg_NrMaxRules(TagType_config_pkg_NrMaxRules),
		.DataType_WIDTH(WIDTH),
		.NumIn(NUM_OPGROUPS),
		.AxiVldRdy(1'b1)
	) i_arbiter(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(flush_i),
		.rr_i(sv2v_uu_i_arbiter_ext_rr_i_0),
		.req_i(opgrp_out_valid),
		.gnt_o(opgrp_out_ready),
		.data_i(opgrp_outputs),
		.gnt_i(out_ready_i),
		.req_o(out_valid_o),
		.data_o(arbiter_output),
		.idx_o()
	);
	// Trace: core/cvfpu/src/fpnew_top.sv:179:3
	assign result_o = arbiter_output[WIDTH + (TagType_CVA6Cfg[8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 4)-:((WIDTH + (TagType_CVA6Cfg[8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 4)) >= (5 + (TagType_CVA6Cfg[8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0)) ? ((WIDTH + (TagType_CVA6Cfg[8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 4)) - (5 + (TagType_CVA6Cfg[8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0))) + 1 : ((5 + (TagType_CVA6Cfg[8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0)) - (WIDTH + (TagType_CVA6Cfg[8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 4))) + 1)];
	// Trace: core/cvfpu/src/fpnew_top.sv:180:3
	assign status_o = arbiter_output[TagType_CVA6Cfg[8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 4-:((TagType_CVA6Cfg[8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 4) >= (TagType_CVA6Cfg[8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0) ? ((TagType_CVA6Cfg[8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 4) - (TagType_CVA6Cfg[8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0)) + 1 : ((TagType_CVA6Cfg[8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0) - (TagType_CVA6Cfg[8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 4)) + 1)];
	// Trace: core/cvfpu/src/fpnew_top.sv:181:3
	assign tag_o = arbiter_output[TagType_CVA6Cfg[8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1-:TagType_CVA6Cfg[8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_config_pkg_NrMaxRules * 64) + ((TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]];
	// Trace: core/cvfpu/src/fpnew_top.sv:183:3
	assign busy_o = |opgrp_busy;
	initial _sv2v_0 = 0;
endmodule
