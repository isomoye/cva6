// removed module with interface ports: axi_join_intf
