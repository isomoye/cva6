module id_stage_1271B_A4180 (
	clk_i,
	rst_ni,
	flush_i,
	debug_req_i,
	fetch_entry_i,
	fetch_entry_valid_i,
	fetch_entry_ready_o,
	issue_entry_o,
	orig_instr_o,
	issue_entry_valid_o,
	is_ctrl_flow_o,
	issue_instr_ack_i,
	rvfi_is_compressed_o,
	priv_lvl_i,
	v_i,
	fs_i,
	vfs_i,
	frm_i,
	vs_i,
	irq_i,
	irq_ctrl_i,
	debug_mode_i,
	tvm_i,
	tw_i,
	vtw_i,
	tsr_i,
	hu_i,
	hart_id_i,
	compressed_ready_i,
	compressed_resp_i,
	compressed_valid_o,
	compressed_req_o
);
	// removed localparam type branchpredict_sbe_t_CVA6Cfg_type
	parameter [17102:0] branchpredict_sbe_t_CVA6Cfg = 0;
	// removed localparam type exception_t_CVA6Cfg_type
	parameter [17102:0] exception_t_CVA6Cfg = 0;
	// removed localparam type fetch_entry_t_CVA6Cfg_type
	parameter [17102:0] fetch_entry_t_CVA6Cfg = 0;
	// removed localparam type interrupts_t_CVA6Cfg_type
	parameter [17102:0] interrupts_t_CVA6Cfg = 0;
	// removed localparam type irq_ctrl_t_CVA6Cfg_type
	parameter [17102:0] irq_ctrl_t_CVA6Cfg = 0;
	// removed localparam type scoreboard_entry_t_CVA6Cfg_type
	parameter [17102:0] scoreboard_entry_t_CVA6Cfg = 0;
	// removed localparam type x_compressed_req_t_x_compressed_req_t_CVA6Cfg_type
	parameter [17102:0] x_compressed_req_t_x_compressed_req_t_CVA6Cfg = 0;
	reg _sv2v_0;
	// Trace: core/id_stage.sv:17:15
	localparam config_pkg_NrMaxRules = 16;
	// removed localparam type config_pkg_cache_type_t
	// removed localparam type config_pkg_noc_type_e
	// removed localparam type config_pkg_vm_mode_t
	// removed localparam type config_pkg_cva6_cfg_t
	localparam [17102:0] config_pkg_cva6_cfg_empty = 17103'd0;
	parameter [17102:0] CVA6Cfg = config_pkg_cva6_cfg_empty;
	// Trace: core/id_stage.sv:18:20
	// removed localparam type branchpredict_sbe_t
	// Trace: core/id_stage.sv:19:20
	// removed localparam type exception_t
	// Trace: core/id_stage.sv:20:20
	// removed localparam type fetch_entry_t
	// Trace: core/id_stage.sv:21:20
	// removed localparam type irq_ctrl_t
	// Trace: core/id_stage.sv:22:20
	// removed localparam type scoreboard_entry_t
	// Trace: core/id_stage.sv:23:20
	// removed localparam type interrupts_t
	// Trace: core/id_stage.sv:24:15
	parameter [(((((((((interrupts_t_CVA6Cfg[17102-:32] + interrupts_t_CVA6Cfg[17102-:32]) + interrupts_t_CVA6Cfg[17102-:32]) + interrupts_t_CVA6Cfg[17102-:32]) + interrupts_t_CVA6Cfg[17102-:32]) + interrupts_t_CVA6Cfg[17102-:32]) + interrupts_t_CVA6Cfg[17102-:32]) + interrupts_t_CVA6Cfg[17102-:32]) + interrupts_t_CVA6Cfg[17102-:32]) + interrupts_t_CVA6Cfg[17102-:32]) - 1:0] INTERRUPTS = 1'sb0;
	// Trace: core/id_stage.sv:25:20
	// removed localparam type x_compressed_req_t
	// Trace: core/id_stage.sv:26:20
	// removed localparam type x_compressed_resp_t
	// Trace: core/id_stage.sv:29:5
	input wire clk_i;
	// Trace: core/id_stage.sv:31:5
	input wire rst_ni;
	// Trace: core/id_stage.sv:33:5
	input wire flush_i;
	// Trace: core/id_stage.sv:35:5
	input wire debug_req_i;
	// Trace: core/id_stage.sv:37:5
	input wire [(CVA6Cfg[16841-:32] * (((fetch_entry_t_CVA6Cfg[17070-:32] + 32) + (3 + fetch_entry_t_CVA6Cfg[17070-:32])) + ((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33)))) - 1:0] fetch_entry_i;
	// Trace: core/id_stage.sv:39:5
	input wire [CVA6Cfg[16841-:32] - 1:0] fetch_entry_valid_i;
	// Trace: core/id_stage.sv:41:5
	output reg [CVA6Cfg[16841-:32] - 1:0] fetch_entry_ready_o;
	// Trace: core/id_stage.sv:43:5
	output wire [((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (CVA6Cfg[16841-:32] * (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5)) - 1 : (CVA6Cfg[16841-:32] * (1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 3)):((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 0 : ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)] issue_entry_o;
	// Trace: core/id_stage.sv:45:5
	output wire [(CVA6Cfg[16841-:32] * 32) - 1:0] orig_instr_o;
	// Trace: core/id_stage.sv:47:5
	output wire [CVA6Cfg[16841-:32] - 1:0] issue_entry_valid_o;
	// Trace: core/id_stage.sv:49:5
	output wire [CVA6Cfg[16841-:32] - 1:0] is_ctrl_flow_o;
	// Trace: core/id_stage.sv:51:5
	input wire [CVA6Cfg[16841-:32] - 1:0] issue_instr_ack_i;
	// Trace: core/id_stage.sv:53:5
	output wire [CVA6Cfg[16841-:32] - 1:0] rvfi_is_compressed_o;
	// Trace: core/id_stage.sv:55:5
	// removed localparam type riscv_priv_lvl_t
	input wire [1:0] priv_lvl_i;
	// Trace: core/id_stage.sv:57:5
	input wire v_i;
	// Trace: core/id_stage.sv:59:5
	// removed localparam type riscv_xs_t
	input wire [1:0] fs_i;
	// Trace: core/id_stage.sv:61:5
	input wire [1:0] vfs_i;
	// Trace: core/id_stage.sv:63:5
	input wire [2:0] frm_i;
	// Trace: core/id_stage.sv:65:5
	input wire [1:0] vs_i;
	// Trace: core/id_stage.sv:67:5
	input wire [1:0] irq_i;
	// Trace: core/id_stage.sv:69:5
	input wire [(((irq_ctrl_t_CVA6Cfg[17102-:32] + irq_ctrl_t_CVA6Cfg[17102-:32]) + irq_ctrl_t_CVA6Cfg[17102-:32]) + irq_ctrl_t_CVA6Cfg[17102-:32]) + 1:0] irq_ctrl_i;
	// Trace: core/id_stage.sv:71:5
	input wire debug_mode_i;
	// Trace: core/id_stage.sv:73:5
	input wire tvm_i;
	// Trace: core/id_stage.sv:75:5
	input wire tw_i;
	// Trace: core/id_stage.sv:77:5
	input wire vtw_i;
	// Trace: core/id_stage.sv:79:5
	input wire tsr_i;
	// Trace: core/id_stage.sv:81:5
	input wire hu_i;
	// Trace: core/id_stage.sv:83:5
	input wire [CVA6Cfg[17102-:32] - 1:0] hart_id_i;
	// Trace: core/id_stage.sv:84:5
	input wire compressed_ready_i;
	// Trace: core/id_stage.sv:85:5
	input wire [32:0] compressed_resp_i;
	// Trace: core/id_stage.sv:86:5
	output wire compressed_valid_o;
	// Trace: core/id_stage.sv:87:5
	output wire [(16 + x_compressed_req_t_x_compressed_req_t_CVA6Cfg[127-:32]) - 1:0] compressed_req_o;
	// Trace: core/id_stage.sv:90:3
	// removed localparam type issue_struct_t
	// Trace: core/id_stage.sv:96:3
	reg [(((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) >= 0 ? (CVA6Cfg[16841-:32] * ((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 33)) - 1 : (CVA6Cfg[16841-:32] * (1 - ((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32))) + ((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 31)):(((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) >= 0 ? 0 : (1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32)] issue_n;
	reg [(((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) >= 0 ? (CVA6Cfg[16841-:32] * ((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 33)) - 1 : (CVA6Cfg[16841-:32] * (1 - ((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32))) + ((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 31)):(((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) >= 0 ? 0 : (1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32)] issue_q;
	// Trace: core/id_stage.sv:98:3
	wire [CVA6Cfg[16841-:32] - 1:0] is_control_flow_instr;
	// Trace: core/id_stage.sv:99:3
	wire [((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (CVA6Cfg[16841-:32] * (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5)) - 1 : (CVA6Cfg[16841-:32] * (1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 3)):((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 0 : ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)] decoded_instruction;
	// Trace: core/id_stage.sv:100:3
	wire [(CVA6Cfg[16841-:32] * 32) - 1:0] orig_instr;
	// Trace: core/id_stage.sv:102:3
	wire [CVA6Cfg[16841-:32] - 1:0] is_illegal;
	// Trace: core/id_stage.sv:103:3
	wire [CVA6Cfg[16841-:32] - 1:0] is_illegal_cmp;
	// Trace: core/id_stage.sv:104:3
	wire [CVA6Cfg[16841-:32] - 1:0] is_illegal_cvxif;
	// Trace: core/id_stage.sv:105:3
	wire [(CVA6Cfg[16841-:32] * 32) - 1:0] instruction;
	// Trace: core/id_stage.sv:106:3
	wire [(CVA6Cfg[16841-:32] * 32) - 1:0] compressed_instr;
	// Trace: core/id_stage.sv:107:3
	wire [(CVA6Cfg[16841-:32] * 32) - 1:0] instruction_cvxif;
	// Trace: core/id_stage.sv:108:3
	wire [CVA6Cfg[16841-:32] - 1:0] is_compressed;
	// Trace: core/id_stage.sv:109:3
	wire [CVA6Cfg[16841-:32] - 1:0] is_compressed_cmp;
	// Trace: core/id_stage.sv:110:3
	wire [CVA6Cfg[16841-:32] - 1:0] is_compressed_cvxif;
	// Trace: core/id_stage.sv:112:3
	wire [CVA6Cfg[16841-:32] - 1:0] is_macro_instr_i;
	// Trace: core/id_stage.sv:113:3
	wire stall_instr_fetch;
	// Trace: core/id_stage.sv:114:3
	wire stall_macro_deco;
	// Trace: core/id_stage.sv:115:3
	wire is_last_macro_instr_o;
	// Trace: core/id_stage.sv:116:3
	wire is_double_rd_macro_instr_o;
	// Trace: core/id_stage.sv:118:3
	generate
		if (CVA6Cfg[16544]) begin : genblk1
			genvar _gv_i_20;
			for (_gv_i_20 = 0; _gv_i_20 < CVA6Cfg[16841-:32]; _gv_i_20 = _gv_i_20 + 1) begin : genblk1
				localparam i = _gv_i_20;
				// Trace: core/id_stage.sv:123:7
				compressed_decoder #(.CVA6Cfg(CVA6Cfg)) compressed_decoder_i(
					.instr_i(fetch_entry_i[(i * (((fetch_entry_t_CVA6Cfg[17070-:32] + 32) + (3 + fetch_entry_t_CVA6Cfg[17070-:32])) + ((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33)))) + (32 + ((3 + fetch_entry_t_CVA6Cfg[17070-:32]) + (((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33)) - 1)))-:((32 + ((3 + fetch_entry_t_CVA6Cfg[17070-:32]) + (((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33)) - 1))) >= ((3 + fetch_entry_t_CVA6Cfg[17070-:32]) + (((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33)) + 0)) ? ((32 + ((3 + fetch_entry_t_CVA6Cfg[17070-:32]) + (((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33)) - 1))) - ((3 + fetch_entry_t_CVA6Cfg[17070-:32]) + (((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33)) + 0))) + 1 : (((3 + fetch_entry_t_CVA6Cfg[17070-:32]) + (((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33)) + 0)) - (32 + ((3 + fetch_entry_t_CVA6Cfg[17070-:32]) + (((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33)) - 1)))) + 1)]),
					.instr_o(compressed_instr[i * 32+:32]),
					.illegal_instr_o(is_illegal[i]),
					.is_compressed_o(is_compressed[i]),
					.is_macro_instr_o(is_macro_instr_i[i])
				);
			end
			if (CVA6Cfg[16541]) begin : genblk2
				// Trace: core/id_stage.sv:135:7
				macro_decoder #(.CVA6Cfg(CVA6Cfg)) macro_decoder_i(
					.instr_i(compressed_instr[0+:32]),
					.is_macro_instr_i(is_macro_instr_i[0]),
					.clk_i(clk_i),
					.rst_ni(rst_ni),
					.instr_o(instruction_cvxif[0+:32]),
					.illegal_instr_i(is_illegal[0]),
					.is_compressed_i(is_compressed[0]),
					.issue_ack_i(issue_instr_ack_i[0]),
					.illegal_instr_o(is_illegal_cvxif[0]),
					.is_compressed_o(is_compressed_cvxif[0]),
					.fetch_stall_o(stall_macro_deco),
					.is_last_macro_instr_o(is_last_macro_instr_o),
					.is_double_rd_macro_instr_o(is_double_rd_macro_instr_o)
				);
				if (CVA6Cfg[16874]) begin : genblk1
					// Trace: core/id_stage.sv:153:9
					assign instruction_cvxif[(CVA6Cfg[16841-:32] - 1) * 32+:32] = 1'sb0;
					// Trace: core/id_stage.sv:154:9
					assign is_illegal_cvxif[CVA6Cfg[16841-:32] - 1] = 1'sb0;
					// Trace: core/id_stage.sv:155:9
					assign is_compressed_cvxif[CVA6Cfg[16841-:32] - 1] = 1'sb0;
				end
				// Trace: core/id_stage.sv:157:7
				cvxif_compressed_if_driver_4B483_D0D6F #(
					.x_compressed_req_t_x_compressed_req_t_x_compressed_req_t_CVA6Cfg(x_compressed_req_t_x_compressed_req_t_CVA6Cfg),
					.CVA6Cfg(CVA6Cfg)
				) i_cvxif_compressed_if_driver_i(
					.clk_i(clk_i),
					.rst_ni(rst_ni),
					.hart_id_i(hart_id_i),
					.is_compressed_i(is_compressed_cvxif),
					.is_illegal_i(is_illegal_cvxif),
					.instruction_i(instruction_cvxif),
					.is_compressed_o(is_compressed_cmp),
					.is_illegal_o(is_illegal_cmp),
					.instruction_o(instruction),
					.stall_i(stall_macro_deco),
					.stall_o(stall_instr_fetch),
					.compressed_ready_i(compressed_ready_i),
					.compressed_resp_i(compressed_resp_i),
					.compressed_valid_o(compressed_valid_o),
					.compressed_req_o(compressed_req_o)
				);
			end
			else begin : genblk2
				// Trace: core/id_stage.sv:179:7
				cvxif_compressed_if_driver_4B483_D0D6F #(
					.x_compressed_req_t_x_compressed_req_t_x_compressed_req_t_CVA6Cfg(x_compressed_req_t_x_compressed_req_t_CVA6Cfg),
					.CVA6Cfg(CVA6Cfg)
				) i_cvxif_compressed_if_driver_i(
					.clk_i(clk_i),
					.rst_ni(rst_ni),
					.hart_id_i(hart_id_i),
					.is_compressed_i(is_compressed),
					.is_illegal_i(is_illegal),
					.instruction_i(compressed_instr),
					.is_compressed_o(is_compressed_cmp),
					.is_illegal_o(is_illegal_cmp),
					.instruction_o(instruction),
					.stall_i(1'b0),
					.stall_o(stall_instr_fetch),
					.compressed_ready_i(compressed_ready_i),
					.compressed_resp_i(compressed_resp_i),
					.compressed_valid_o(compressed_valid_o),
					.compressed_req_o(compressed_req_o)
				);
				// Trace: core/id_stage.sv:200:7
				assign is_last_macro_instr_o = 1'sb0;
				// Trace: core/id_stage.sv:201:7
				assign is_double_rd_macro_instr_o = 1'sb0;
			end
		end
		else begin : genblk1
			genvar _gv_i_21;
			for (_gv_i_21 = 0; _gv_i_21 < CVA6Cfg[16841-:32]; _gv_i_21 = _gv_i_21 + 1) begin : genblk1
				localparam i = _gv_i_21;
				// Trace: core/id_stage.sv:205:7
				assign instruction[i * 32+:32] = fetch_entry_i[(i * (((fetch_entry_t_CVA6Cfg[17070-:32] + 32) + (3 + fetch_entry_t_CVA6Cfg[17070-:32])) + ((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33)))) + (32 + ((3 + fetch_entry_t_CVA6Cfg[17070-:32]) + (((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33)) - 1)))-:((32 + ((3 + fetch_entry_t_CVA6Cfg[17070-:32]) + (((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33)) - 1))) >= ((3 + fetch_entry_t_CVA6Cfg[17070-:32]) + (((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33)) + 0)) ? ((32 + ((3 + fetch_entry_t_CVA6Cfg[17070-:32]) + (((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33)) - 1))) - ((3 + fetch_entry_t_CVA6Cfg[17070-:32]) + (((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33)) + 0))) + 1 : (((3 + fetch_entry_t_CVA6Cfg[17070-:32]) + (((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33)) + 0)) - (32 + ((3 + fetch_entry_t_CVA6Cfg[17070-:32]) + (((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33)) - 1)))) + 1)];
			end
			// Trace: core/id_stage.sv:207:5
			assign is_illegal_cmp = 1'sb0;
			// Trace: core/id_stage.sv:208:5
			assign is_compressed_cmp = 1'sb0;
			// Trace: core/id_stage.sv:209:5
			assign is_macro_instr_i = 1'sb0;
			// Trace: core/id_stage.sv:210:5
			assign is_last_macro_instr_o = 1'sb0;
			// Trace: core/id_stage.sv:211:5
			assign is_double_rd_macro_instr_o = 1'sb0;
			if (CVA6Cfg[16539]) begin : genblk2
				// Trace: core/id_stage.sv:213:7
				assign compressed_valid_o = 1'sb0;
				// Trace: core/id_stage.sv:214:7
				assign compressed_req_o[x_compressed_req_t_x_compressed_req_t_CVA6Cfg[127-:32] + 15-:((x_compressed_req_t_x_compressed_req_t_CVA6Cfg[127-:32] + 15) >= (x_compressed_req_t_x_compressed_req_t_CVA6Cfg[127-:32] + 0) ? ((x_compressed_req_t_x_compressed_req_t_CVA6Cfg[127-:32] + 15) - (x_compressed_req_t_x_compressed_req_t_CVA6Cfg[127-:32] + 0)) + 1 : ((x_compressed_req_t_x_compressed_req_t_CVA6Cfg[127-:32] + 0) - (x_compressed_req_t_x_compressed_req_t_CVA6Cfg[127-:32] + 15)) + 1)] = 1'sb0;
				// Trace: core/id_stage.sv:215:7
				assign compressed_req_o[x_compressed_req_t_x_compressed_req_t_CVA6Cfg[127-:32] - 1-:x_compressed_req_t_x_compressed_req_t_CVA6Cfg[127-:32]] = hart_id_i;
			end
		end
	endgenerate
	// Trace: core/id_stage.sv:219:3
	assign rvfi_is_compressed_o = is_compressed_cmp;
	// Trace: core/id_stage.sv:223:3
	genvar _gv_i_22;
	generate
		for (_gv_i_22 = 0; _gv_i_22 < CVA6Cfg[16841-:32]; _gv_i_22 = _gv_i_22 + 1) begin : genblk2
			localparam i = _gv_i_22;
			// Trace: core/id_stage.sv:224:5
			decoder_90836_06260 #(
				.branchpredict_sbe_t_branchpredict_sbe_t_CVA6Cfg(branchpredict_sbe_t_CVA6Cfg),
				.exception_t_exception_t_CVA6Cfg(exception_t_CVA6Cfg),
				.interrupts_t_interrupts_t_CVA6Cfg(interrupts_t_CVA6Cfg),
				.irq_ctrl_t_irq_ctrl_t_CVA6Cfg(irq_ctrl_t_CVA6Cfg),
				.scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg(scoreboard_entry_t_CVA6Cfg),
				.CVA6Cfg(CVA6Cfg),
				.INTERRUPTS(INTERRUPTS)
			) decoder_i(
				.debug_req_i(debug_req_i),
				.irq_ctrl_i(irq_ctrl_i),
				.irq_i(irq_i),
				.pc_i(fetch_entry_i[(i * (((fetch_entry_t_CVA6Cfg[17070-:32] + 32) + (3 + fetch_entry_t_CVA6Cfg[17070-:32])) + ((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33)))) + (fetch_entry_t_CVA6Cfg[17070-:32] + (32 + ((3 + fetch_entry_t_CVA6Cfg[17070-:32]) + (((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33)) - 1))))-:((fetch_entry_t_CVA6Cfg[17070-:32] + (32 + ((3 + fetch_entry_t_CVA6Cfg[17070-:32]) + (((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33)) - 1)))) >= (32 + ((3 + fetch_entry_t_CVA6Cfg[17070-:32]) + (((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33)) + 0))) ? ((fetch_entry_t_CVA6Cfg[17070-:32] + (32 + ((3 + fetch_entry_t_CVA6Cfg[17070-:32]) + (((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33)) - 1)))) - (32 + ((3 + fetch_entry_t_CVA6Cfg[17070-:32]) + (((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33)) + 0)))) + 1 : ((32 + ((3 + fetch_entry_t_CVA6Cfg[17070-:32]) + (((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33)) + 0))) - (fetch_entry_t_CVA6Cfg[17070-:32] + (32 + ((3 + fetch_entry_t_CVA6Cfg[17070-:32]) + (((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33)) - 1))))) + 1)]),
				.is_compressed_i(is_compressed_cmp[i]),
				.is_macro_instr_i(is_macro_instr_i[i]),
				.is_last_macro_instr_i(is_last_macro_instr_o),
				.is_double_rd_macro_instr_i(is_double_rd_macro_instr_o),
				.is_illegal_i(is_illegal_cmp[i]),
				.instruction_i(instruction[i * 32+:32]),
				.compressed_instr_i(fetch_entry_i[(i * (((fetch_entry_t_CVA6Cfg[17070-:32] + 32) + (3 + fetch_entry_t_CVA6Cfg[17070-:32])) + ((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33)))) + (((32 + ((3 + fetch_entry_t_CVA6Cfg[17070-:32]) + (((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33)) - 1))) - 16) >= ((32 + ((3 + fetch_entry_t_CVA6Cfg[17070-:32]) + (((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33)) - 1))) - 31) ? (32 + ((3 + fetch_entry_t_CVA6Cfg[17070-:32]) + (((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33)) - 1))) - 16 : (((32 + ((3 + fetch_entry_t_CVA6Cfg[17070-:32]) + (((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33)) - 1))) - 16) + (((32 + ((3 + fetch_entry_t_CVA6Cfg[17070-:32]) + (((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33)) - 1))) - 16) >= ((32 + ((3 + fetch_entry_t_CVA6Cfg[17070-:32]) + (((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33)) - 1))) - 31) ? (((32 + ((3 + fetch_entry_t_CVA6Cfg[17070-:32]) + (((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33)) - 1))) - 16) - ((32 + ((3 + fetch_entry_t_CVA6Cfg[17070-:32]) + (((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33)) - 1))) - 31)) + 1 : (((32 + ((3 + fetch_entry_t_CVA6Cfg[17070-:32]) + (((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33)) - 1))) - 31) - ((32 + ((3 + fetch_entry_t_CVA6Cfg[17070-:32]) + (((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33)) - 1))) - 16)) + 1)) - 1)-:(((32 + ((3 + fetch_entry_t_CVA6Cfg[17070-:32]) + (((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33)) - 1))) - 16) >= ((32 + ((3 + fetch_entry_t_CVA6Cfg[17070-:32]) + (((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33)) - 1))) - 31) ? (((32 + ((3 + fetch_entry_t_CVA6Cfg[17070-:32]) + (((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33)) - 1))) - 16) - ((32 + ((3 + fetch_entry_t_CVA6Cfg[17070-:32]) + (((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33)) - 1))) - 31)) + 1 : (((32 + ((3 + fetch_entry_t_CVA6Cfg[17070-:32]) + (((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33)) - 1))) - 31) - ((32 + ((3 + fetch_entry_t_CVA6Cfg[17070-:32]) + (((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33)) - 1))) - 16)) + 1)]),
				.branch_predict_i(fetch_entry_i[(i * (((fetch_entry_t_CVA6Cfg[17070-:32] + 32) + (3 + fetch_entry_t_CVA6Cfg[17070-:32])) + ((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33)))) + ((3 + fetch_entry_t_CVA6Cfg[17070-:32]) + (((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33)) - 1))-:(((3 + fetch_entry_t_CVA6Cfg[17070-:32]) + (((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33)) - 1)) >= (((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33)) + 0) ? (((3 + fetch_entry_t_CVA6Cfg[17070-:32]) + (((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33)) - 1)) - (((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33)) + 0)) + 1 : ((((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33)) + 0) - ((3 + fetch_entry_t_CVA6Cfg[17070-:32]) + (((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33)) - 1))) + 1)]),
				.ex_i(fetch_entry_i[(i * (((fetch_entry_t_CVA6Cfg[17070-:32] + 32) + (3 + fetch_entry_t_CVA6Cfg[17070-:32])) + ((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33)))) + (((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33)) - 1)-:((((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((fetch_entry_t_CVA6Cfg[17102-:32] + fetch_entry_t_CVA6Cfg[17102-:32]) + fetch_entry_t_CVA6Cfg[17006-:32]) + 33))]),
				.priv_lvl_i(priv_lvl_i),
				.v_i(v_i),
				.debug_mode_i(debug_mode_i),
				.fs_i(fs_i),
				.vfs_i(vfs_i),
				.frm_i(frm_i),
				.vs_i(vs_i),
				.tvm_i(tvm_i),
				.tw_i(tw_i),
				.vtw_i(vtw_i),
				.tsr_i(tsr_i),
				.hu_i(hu_i),
				.instruction_o(decoded_instruction[((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 0 : ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) + (i * ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))+:((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))]),
				.orig_instr_o(orig_instr[i * 32+:32]),
				.is_control_flow_instr_o(is_control_flow_instr[i])
			);
		end
	endgenerate
	// Trace: core/id_stage.sv:267:3
	genvar _gv_i_23;
	generate
		for (_gv_i_23 = 0; _gv_i_23 < CVA6Cfg[16841-:32]; _gv_i_23 = _gv_i_23 + 1) begin : genblk3
			localparam i = _gv_i_23;
			// Trace: core/id_stage.sv:268:5
			assign issue_entry_o[((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 0 : ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) + (i * ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))+:((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))] = issue_q[(((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) >= 0 ? (i * (((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) >= 0 ? (1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 33 : 1 - ((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32))) + (((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) >= 0 ? ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 32 : ((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) - (((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 32)) : (((i * (((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) >= 0 ? (1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 33 : 1 - ((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32))) + (((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) >= 0 ? ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 32 : ((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) - (((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 32))) + ((((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 32) >= 33 ? ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 0 : 34 - (((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 32))) - 1)-:((((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 32) >= 33 ? ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 0 : 34 - (((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 32))];
			// Trace: core/id_stage.sv:269:5
			assign issue_entry_valid_o[i] = issue_q[(i * (((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) >= 0 ? (1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 33 : 1 - ((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32))) + (((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) >= 0 ? 1 + (((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 32) : ((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) - (1 + (((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 32)))];
			// Trace: core/id_stage.sv:270:5
			assign is_ctrl_flow_o[i] = issue_q[(i * (((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) >= 0 ? (1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 33 : 1 - ((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32))) + (((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) >= 0 ? 0 : (1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32)];
			// Trace: core/id_stage.sv:271:5
			assign orig_instr_o[i * 32+:32] = issue_q[(((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) >= 0 ? (i * (((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) >= 0 ? (1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 33 : 1 - ((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32))) + (((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) >= 0 ? 32 : (1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 0) : ((i * (((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) >= 0 ? (1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 33 : 1 - ((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32))) + (((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) >= 0 ? 32 : (1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 0)) + 31)-:32];
		end
	endgenerate
	// Trace: core/id_stage.sv:274:3
	generate
		if (CVA6Cfg[16874]) begin : genblk4
			// Trace: core/id_stage.sv:275:5
			always @(*) begin
				if (_sv2v_0)
					;
				// Trace: core/id_stage.sv:276:7
				issue_n = issue_q;
				// Trace: core/id_stage.sv:277:7
				fetch_entry_ready_o = 1'sb0;
				// Trace: core/id_stage.sv:280:7
				if (issue_instr_ack_i[0])
					// Trace: core/id_stage.sv:281:9
					issue_n[0 + (((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) >= 0 ? 1 + (((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 32) : ((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) - (1 + (((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 32)))] = 1'b0;
				if (issue_instr_ack_i[1])
					// Trace: core/id_stage.sv:284:9
					issue_n[(((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) >= 0 ? (1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 33 : 1 - ((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32)) + (((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) >= 0 ? 1 + (((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 32) : ((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) - (1 + (((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 32)))] = 1'b0;
				if (!issue_n[0 + (((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) >= 0 ? 1 + (((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 32) : ((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) - (1 + (((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 32)))]) begin
					begin
						// Trace: core/id_stage.sv:288:9
						if (issue_n[(((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) >= 0 ? (1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 33 : 1 - ((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32)) + (((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) >= 0 ? 1 + (((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 32) : ((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) - (1 + (((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 32)))]) begin
							// Trace: core/id_stage.sv:289:11
							issue_n[(((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) >= 0 ? 0 : (1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) + 0+:(((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) >= 0 ? (1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 33 : 1 - ((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32))] = issue_n[(((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) >= 0 ? 0 : (1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) + (((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) >= 0 ? (1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 33 : 1 - ((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32))+:(((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) >= 0 ? (1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 33 : 1 - ((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32))];
							// Trace: core/id_stage.sv:290:11
							issue_n[(((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) >= 0 ? (1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 33 : 1 - ((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32)) + (((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) >= 0 ? 1 + (((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 32) : ((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) - (1 + (((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 32)))] = 1'b0;
						end
						else if (fetch_entry_valid_i[0]) begin
							// Trace: core/id_stage.sv:292:11
							fetch_entry_ready_o[0] = 1'b1;
							// Trace: core/id_stage.sv:293:11
							issue_n[(((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) >= 0 ? 0 : (1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) + 0+:(((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) >= 0 ? (1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 33 : 1 - ((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32))] = {1'b1, decoded_instruction[((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 0 : ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) + 0+:((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))], orig_instr[0+:32], is_control_flow_instr[0]};
						end
					end
				end
				if (!issue_n[(((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) >= 0 ? (1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 33 : 1 - ((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32)) + (((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) >= 0 ? 1 + (((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 32) : ((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) - (1 + (((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 32)))]) begin
					begin
						// Trace: core/id_stage.sv:298:9
						if (fetch_entry_ready_o[0]) begin
							begin
								// Trace: core/id_stage.sv:299:11
								if (fetch_entry_valid_i[1]) begin
									// Trace: core/id_stage.sv:300:13
									fetch_entry_ready_o[1] = 1'b1;
									// Trace: core/id_stage.sv:301:13
									issue_n[(((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) >= 0 ? 0 : (1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) + (((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) >= 0 ? (1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 33 : 1 - ((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32))+:(((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) >= 0 ? (1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 33 : 1 - ((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32))] = {1'b1, decoded_instruction[((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 0 : ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))+:((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))], orig_instr[32+:32], is_control_flow_instr[1]};
								end
							end
						end
						else if (fetch_entry_valid_i[0]) begin
							// Trace: core/id_stage.sv:304:11
							fetch_entry_ready_o[0] = 1'b1;
							// Trace: core/id_stage.sv:305:11
							issue_n[(((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) >= 0 ? 0 : (1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) + (((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) >= 0 ? (1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 33 : 1 - ((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32))+:(((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) >= 0 ? (1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 33 : 1 - ((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32))] = {1'b1, decoded_instruction[((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 0 : ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) + 0+:((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))], orig_instr[0+:32], is_control_flow_instr[0]};
						end
					end
				end
				if (flush_i) begin
					// Trace: core/id_stage.sv:310:9
					issue_n[0 + (((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) >= 0 ? 1 + (((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 32) : ((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) - (1 + (((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 32)))] = 1'b0;
					// Trace: core/id_stage.sv:311:9
					issue_n[(((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) >= 0 ? (1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 33 : 1 - ((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32)) + (((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) >= 0 ? 1 + (((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 32) : ((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) - (1 + (((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 32)))] = 1'b0;
				end
			end
		end
		else begin : genblk4
			// Trace: core/id_stage.sv:315:5
			always @(*) begin
				if (_sv2v_0)
					;
				// Trace: core/id_stage.sv:316:7
				issue_n = issue_q;
				// Trace: core/id_stage.sv:317:7
				fetch_entry_ready_o = 1'sb0;
				// Trace: core/id_stage.sv:320:7
				if (issue_instr_ack_i[0])
					// Trace: core/id_stage.sv:320:33
					issue_n[0 + (((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) >= 0 ? 1 + (((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 32) : ((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) - (1 + (((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 32)))] = 1'b0;
				if ((!issue_q[0 + (((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) >= 0 ? 1 + (((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 32) : ((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) - (1 + (((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 32)))] || issue_instr_ack_i[0]) && fetch_entry_valid_i[0]) begin
					// Trace: core/id_stage.sv:326:9
					if (stall_instr_fetch)
						// Trace: core/id_stage.sv:327:11
						fetch_entry_ready_o[0] = 1'b0;
					else
						// Trace: core/id_stage.sv:329:11
						fetch_entry_ready_o[0] = 1'b1;
					// Trace: core/id_stage.sv:331:9
					issue_n[(((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) >= 0 ? 0 : (1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) + 0+:(((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) >= 0 ? (1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 33 : 1 - ((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32))] = {1'b1, decoded_instruction[((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 0 : ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) + 0+:((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))], orig_instr[0+:32], is_control_flow_instr[0]};
				end
				if (flush_i)
					// Trace: core/id_stage.sv:335:20
					issue_n[0 + (((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) >= 0 ? 1 + (((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 32) : ((1 + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + 32) - (1 + (((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 32)))] = 1'b0;
			end
		end
	endgenerate
	// Trace: core/id_stage.sv:341:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: core/id_stage.sv:342:5
		if (~rst_ni)
			// Trace: core/id_stage.sv:343:7
			issue_q <= 1'sb0;
		else
			// Trace: core/id_stage.sv:345:7
			issue_q <= issue_n;
	initial _sv2v_0 = 0;
endmodule
