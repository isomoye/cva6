module ras_091E3_171B5 (
	clk_i,
	rst_ni,
	flush_bp_i,
	push_i,
	pop_i,
	data_i,
	data_o
);
	// removed localparam type ras_t_CVA6Cfg_type
	// removed localparam type ras_t_config_pkg_NrMaxRules_type
	parameter [17102:0] ras_t_CVA6Cfg = 0;
	parameter signed [31:0] ras_t_config_pkg_NrMaxRules = 0;
	reg _sv2v_0;
	// Trace: core/frontend/ras.sv:18:15
	localparam config_pkg_NrMaxRules = 16;
	// removed localparam type config_pkg_cache_type_t
	// removed localparam type config_pkg_noc_type_e
	// removed localparam type config_pkg_vm_mode_t
	// removed localparam type config_pkg_cva6_cfg_t
	localparam [17102:0] config_pkg_cva6_cfg_empty = 17103'd0;
	parameter [17102:0] CVA6Cfg = config_pkg_cva6_cfg_empty;
	// Trace: core/frontend/ras.sv:19:20
	// removed localparam type ras_t
	// Trace: core/frontend/ras.sv:20:15
	parameter [31:0] DEPTH = 2;
	// Trace: core/frontend/ras.sv:23:5
	input wire clk_i;
	// Trace: core/frontend/ras.sv:25:5
	input wire rst_ni;
	// Trace: core/frontend/ras.sv:27:5
	input wire flush_bp_i;
	// Trace: core/frontend/ras.sv:29:5
	input wire push_i;
	// Trace: core/frontend/ras.sv:31:5
	input wire pop_i;
	// Trace: core/frontend/ras.sv:33:5
	input wire [CVA6Cfg[17070-:32] - 1:0] data_i;
	// Trace: core/frontend/ras.sv:35:5
	output wire [(1 + ras_t_CVA6Cfg[9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) - 1:0] data_o;
	// Trace: core/frontend/ras.sv:38:3
	reg [(DEPTH * (1 + ras_t_CVA6Cfg[9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)])) - 1:0] stack_d;
	reg [(DEPTH * (1 + ras_t_CVA6Cfg[9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)])) - 1:0] stack_q;
	// Trace: core/frontend/ras.sv:40:3
	assign data_o = stack_q[0+:1 + ras_t_CVA6Cfg[9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]];
	// Trace: core/frontend/ras.sv:42:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: core/frontend/ras.sv:43:5
		stack_d = stack_q;
		// Trace: core/frontend/ras.sv:46:5
		if (push_i) begin
			// Trace: core/frontend/ras.sv:47:7
			stack_d[ras_t_CVA6Cfg[9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1-:ras_t_CVA6Cfg[9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]] = data_i;
			// Trace: core/frontend/ras.sv:49:7
			stack_d[0 + (ras_t_CVA6Cfg[9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0)] = 1'b1;
			// Trace: core/frontend/ras.sv:50:7
			stack_d[(1 + ras_t_CVA6Cfg[9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) * (((DEPTH - 1) >= 1 ? DEPTH - 1 : ((DEPTH - 1) + ((DEPTH - 1) >= 1 ? DEPTH - 1 : 3 - DEPTH)) - 1) - (((DEPTH - 1) >= 1 ? DEPTH - 1 : 3 - DEPTH) - 1))+:(1 + ras_t_CVA6Cfg[9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) * ((DEPTH - 1) >= 1 ? DEPTH - 1 : 3 - DEPTH)] = stack_q[(1 + ras_t_CVA6Cfg[9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) * (((DEPTH - 2) >= 0 ? DEPTH - 2 : ((DEPTH - 2) + ((DEPTH - 2) >= 0 ? DEPTH - 1 : 3 - DEPTH)) - 1) - (((DEPTH - 2) >= 0 ? DEPTH - 1 : 3 - DEPTH) - 1))+:(1 + ras_t_CVA6Cfg[9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) * ((DEPTH - 2) >= 0 ? DEPTH - 1 : 3 - DEPTH)];
		end
		if (pop_i) begin
			// Trace: core/frontend/ras.sv:54:7
			stack_d[(1 + ras_t_CVA6Cfg[9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) * (((DEPTH - 2) >= 0 ? DEPTH - 2 : ((DEPTH - 2) + ((DEPTH - 2) >= 0 ? DEPTH - 1 : 3 - DEPTH)) - 1) - (((DEPTH - 2) >= 0 ? DEPTH - 1 : 3 - DEPTH) - 1))+:(1 + ras_t_CVA6Cfg[9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) * ((DEPTH - 2) >= 0 ? DEPTH - 1 : 3 - DEPTH)] = stack_q[(1 + ras_t_CVA6Cfg[9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) * (((DEPTH - 1) >= 1 ? DEPTH - 1 : ((DEPTH - 1) + ((DEPTH - 1) >= 1 ? DEPTH - 1 : 3 - DEPTH)) - 1) - (((DEPTH - 1) >= 1 ? DEPTH - 1 : 3 - DEPTH) - 1))+:(1 + ras_t_CVA6Cfg[9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) * ((DEPTH - 1) >= 1 ? DEPTH - 1 : 3 - DEPTH)];
			// Trace: core/frontend/ras.sv:56:7
			stack_d[((DEPTH - 1) * (1 + ras_t_CVA6Cfg[9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)])) + (ras_t_CVA6Cfg[9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0)] = 1'b0;
			// Trace: core/frontend/ras.sv:57:7
			stack_d[((DEPTH - 1) * (1 + ras_t_CVA6Cfg[9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)])) + (ras_t_CVA6Cfg[9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1)-:ras_t_CVA6Cfg[9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]] = 'b0;
		end
		if (pop_i && push_i) begin
			// Trace: core/frontend/ras.sv:62:7
			stack_d = stack_q;
			// Trace: core/frontend/ras.sv:63:7
			stack_d[ras_t_CVA6Cfg[9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1-:ras_t_CVA6Cfg[9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]] = data_i;
			// Trace: core/frontend/ras.sv:64:7
			stack_d[0 + (ras_t_CVA6Cfg[9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + (32 + ((ras_t_config_pkg_NrMaxRules * 64) + ((ras_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0)] = 1'b1;
		end
		if (flush_bp_i)
			// Trace: core/frontend/ras.sv:68:7
			stack_d = 1'sb0;
	end
	// Trace: core/frontend/ras.sv:72:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: core/frontend/ras.sv:73:5
		if (~rst_ni)
			// Trace: core/frontend/ras.sv:74:7
			stack_q <= 1'sb0;
		else
			// Trace: core/frontend/ras.sv:76:7
			stack_q <= stack_d;
	initial _sv2v_0 = 0;
endmodule
