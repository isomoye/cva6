module fpnew_opgroup_block_D3AB0_1C1E0 (
	clk_i,
	rst_ni,
	operands_i,
	is_boxed_i,
	rnd_mode_i,
	op_i,
	op_mod_i,
	src_fmt_i,
	dst_fmt_i,
	int_fmt_i,
	vectorial_op_i,
	tag_i,
	simd_mask_i,
	in_valid_i,
	in_ready_o,
	flush_i,
	result_o,
	status_o,
	extension_bit_o,
	tag_o,
	out_valid_o,
	out_ready_i,
	busy_o
);
	// removed localparam type TagType_TagType_CVA6Cfg_type
	// removed localparam type TagType_TagType_config_pkg_NrMaxRules_type
	parameter [17102:0] TagType_TagType_CVA6Cfg = 0;
	parameter signed [31:0] TagType_TagType_config_pkg_NrMaxRules = 0;
	reg _sv2v_0;
	// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:17:13
	// removed localparam type fpnew_pkg_opgroup_e
	parameter [1:0] OpGroup = 2'd0;
	// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:19:13
	parameter [31:0] Width = 32;
	// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:20:13
	parameter [0:0] EnableVectors = 1'b1;
	// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:21:13
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	// removed localparam type fpnew_pkg_fmt_logic_t
	parameter [0:4] FpFmtMask = 1'sb1;
	// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:22:13
	localparam [31:0] fpnew_pkg_NUM_INT_FORMATS = 4;
	// removed localparam type fpnew_pkg_ifmt_logic_t
	parameter [0:3] IntFmtMask = 1'sb1;
	// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:23:13
	// removed localparam type fpnew_pkg_fmt_unsigned_t
	parameter [159:0] FmtPipeRegs = {fpnew_pkg_NUM_FP_FORMATS {32'd0}};
	// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:24:13
	// removed localparam type fpnew_pkg_unit_type_t
	// removed localparam type fpnew_pkg_fmt_unit_types_t
	parameter [9:0] FmtUnitTypes = {fpnew_pkg_NUM_FP_FORMATS {2'd1}};
	// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:25:13
	// removed localparam type fpnew_pkg_pipe_config_t
	parameter [1:0] PipeConfig = 2'd0;
	// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:26:41
	// removed localparam type TagType
	// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:27:13
	parameter [31:0] TrueSIMDClass = 0;
	// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:29:14
	localparam [31:0] NUM_FORMATS = fpnew_pkg_NUM_FP_FORMATS;
	// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:30:14
	function automatic [31:0] fpnew_pkg_num_operands;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:379:48
		input reg [1:0] grp;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:380:5
		(* full_case, parallel_case *)
		case (grp)
			2'd0: fpnew_pkg_num_operands = 3;
			2'd1: fpnew_pkg_num_operands = 2;
			2'd2: fpnew_pkg_num_operands = 2;
			2'd3: fpnew_pkg_num_operands = 3;
			default: fpnew_pkg_num_operands = 0;
		endcase
	endfunction
	localparam [31:0] NUM_OPERANDS = fpnew_pkg_num_operands(OpGroup);
	// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:31:14
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	// removed localparam type fpnew_pkg_fp_format_e
	// removed localparam type fpnew_pkg_fp_encoding_t
	localparam [319:0] fpnew_pkg_FP_ENCODINGS = 320'h8000000170000000b00000034000000050000000a00000005000000020000000800000007;
	function automatic [31:0] fpnew_pkg_fp_width;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:304:44
		input reg [2:0] fmt;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:305:5
		fpnew_pkg_fp_width = (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] + fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32]) + 1;
	endfunction
	function automatic signed [31:0] fpnew_pkg_maximum;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:296:34
		input reg signed [31:0] a;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:296:41
		input reg signed [31:0] b;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:297:5
		fpnew_pkg_maximum = (a > b ? a : b);
	endfunction
	function automatic [2:0] sv2v_cast_5D882;
		input reg [2:0] inp;
		sv2v_cast_5D882 = inp;
	endfunction
	function automatic [31:0] fpnew_pkg_max_fp_width;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:309:48
		input reg [0:4] cfg;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:310:5
		reg [31:0] res;
		begin
			res = 0;
			// Trace: core/cvfpu/src/fpnew_pkg.sv:311:5
			begin : sv2v_autoblock_1
				// Trace: core/cvfpu/src/fpnew_pkg.sv:311:10
				reg [31:0] i;
				// Trace: core/cvfpu/src/fpnew_pkg.sv:311:10
				for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
					if (cfg[i])
						// Trace: core/cvfpu/src/fpnew_pkg.sv:313:9
						res = $unsigned(fpnew_pkg_maximum(res, fpnew_pkg_fp_width(sv2v_cast_5D882(i))));
			end
			fpnew_pkg_max_fp_width = res;
		end
	endfunction
	function automatic signed [31:0] fpnew_pkg_minimum;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:292:34
		input reg signed [31:0] a;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:292:41
		input reg signed [31:0] b;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:293:5
		fpnew_pkg_minimum = (a < b ? a : b);
	endfunction
	function automatic [31:0] fpnew_pkg_min_fp_width;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:318:48
		input reg [0:4] cfg;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:319:5
		reg [31:0] res;
		begin
			res = fpnew_pkg_max_fp_width(cfg);
			// Trace: core/cvfpu/src/fpnew_pkg.sv:320:5
			begin : sv2v_autoblock_2
				// Trace: core/cvfpu/src/fpnew_pkg.sv:320:10
				reg [31:0] i;
				// Trace: core/cvfpu/src/fpnew_pkg.sv:320:10
				for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
					if (cfg[i])
						// Trace: core/cvfpu/src/fpnew_pkg.sv:322:9
						res = $unsigned(fpnew_pkg_minimum(res, fpnew_pkg_fp_width(sv2v_cast_5D882(i))));
			end
			fpnew_pkg_min_fp_width = res;
		end
	endfunction
	function automatic [31:0] fpnew_pkg_max_num_lanes;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:395:49
		input reg [31:0] width;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:395:69
		input reg [0:4] cfg;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:395:86
		input reg vec;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:396:5
		fpnew_pkg_max_num_lanes = (vec ? width / fpnew_pkg_min_fp_width(cfg) : 1);
	endfunction
	localparam [31:0] NUM_LANES = fpnew_pkg_max_num_lanes(Width, FpFmtMask, EnableVectors);
	// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:32:27
	// removed localparam type MaskType
	// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:34:3
	input wire clk_i;
	// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:35:3
	input wire rst_ni;
	// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:37:3
	input wire [(NUM_OPERANDS * Width) - 1:0] operands_i;
	// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:38:3
	input wire [(NUM_FORMATS * NUM_OPERANDS) - 1:0] is_boxed_i;
	// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:39:3
	// removed localparam type fpnew_pkg_roundmode_e
	input wire [2:0] rnd_mode_i;
	// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:40:3
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	// removed localparam type fpnew_pkg_operation_e
	input wire [3:0] op_i;
	// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:41:3
	input wire op_mod_i;
	// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:42:3
	input wire [2:0] src_fmt_i;
	// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:43:3
	input wire [2:0] dst_fmt_i;
	// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:44:3
	localparam [31:0] fpnew_pkg_INT_FORMAT_BITS = 2;
	// removed localparam type fpnew_pkg_int_format_e
	input wire [1:0] int_fmt_i;
	// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:45:3
	input wire vectorial_op_i;
	// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:46:3
	input wire [TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1:0] tag_i;
	// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:47:3
	input wire [NUM_LANES - 1:0] simd_mask_i;
	// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:49:3
	input wire in_valid_i;
	// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:50:3
	output wire in_ready_o;
	// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:51:3
	input wire flush_i;
	// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:53:3
	output wire [Width - 1:0] result_o;
	// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:54:3
	// removed localparam type fpnew_pkg_status_t
	output wire [4:0] status_o;
	// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:55:3
	output wire extension_bit_o;
	// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:56:3
	output wire [TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1:0] tag_o;
	// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:58:3
	output wire out_valid_o;
	// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:59:3
	input wire out_ready_i;
	// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:61:3
	output wire busy_o;
	// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:67:3
	// removed localparam type output_t
	// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:75:3
	wire [4:0] fmt_in_ready;
	wire [4:0] fmt_out_valid;
	wire [4:0] fmt_out_ready;
	wire [4:0] fmt_busy;
	// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:76:3
	wire [(5 * ((Width + 6) + TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)])) - 1:0] fmt_outputs;
	// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:81:3
	assign in_ready_o = in_valid_i & fmt_in_ready[dst_fmt_i];
	// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:86:3
	genvar _gv_fmt_9;
	localparam [0:0] fpnew_pkg_DONT_CARE = 1'b1;
	function automatic fpnew_pkg_any_enabled_multi;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:459:46
		input reg [9:0] types;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:459:70
		input reg [0:4] cfg;
		reg [0:1] _sv2v_jump;
		begin
			_sv2v_jump = 2'b00;
			// Trace: core/cvfpu/src/fpnew_pkg.sv:460:5
			begin : sv2v_autoblock_3
				// Trace: core/cvfpu/src/fpnew_pkg.sv:460:10
				reg [31:0] i;
				// Trace: core/cvfpu/src/fpnew_pkg.sv:460:10
				begin : sv2v_autoblock_4
					reg [31:0] _sv2v_value_on_break;
					for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
						if (_sv2v_jump < 2'b10) begin
							_sv2v_jump = 2'b00;
							if (cfg[i] && (types[(4 - i) * 2+:2] == 2'd2)) begin
								fpnew_pkg_any_enabled_multi = 1'b1;
								_sv2v_jump = 2'b11;
							end
							_sv2v_value_on_break = i;
						end
					if (!(_sv2v_jump < 2'b10))
						i = _sv2v_value_on_break;
					if (_sv2v_jump != 2'b11)
						_sv2v_jump = 2'b00;
				end
			end
			if (_sv2v_jump == 2'b00) begin
				fpnew_pkg_any_enabled_multi = 1'b0;
				_sv2v_jump = 2'b11;
			end
		end
	endfunction
	function automatic [2:0] fpnew_pkg_get_first_enabled_multi;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:477:58
		input reg [9:0] types;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:477:82
		input reg [0:4] cfg;
		reg [0:1] _sv2v_jump;
		begin
			_sv2v_jump = 2'b00;
			// Trace: core/cvfpu/src/fpnew_pkg.sv:478:5
			begin : sv2v_autoblock_5
				// Trace: core/cvfpu/src/fpnew_pkg.sv:478:10
				reg [31:0] i;
				// Trace: core/cvfpu/src/fpnew_pkg.sv:478:10
				begin : sv2v_autoblock_6
					reg [31:0] _sv2v_value_on_break;
					for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
						if (_sv2v_jump < 2'b10) begin
							_sv2v_jump = 2'b00;
							if (cfg[i] && (types[(4 - i) * 2+:2] == 2'd2)) begin
								fpnew_pkg_get_first_enabled_multi = sv2v_cast_5D882(i);
								_sv2v_jump = 2'b11;
							end
							_sv2v_value_on_break = i;
						end
					if (!(_sv2v_jump < 2'b10))
						i = _sv2v_value_on_break;
					if (_sv2v_jump != 2'b11)
						_sv2v_jump = 2'b00;
				end
			end
			if (_sv2v_jump == 2'b00) begin
				fpnew_pkg_get_first_enabled_multi = sv2v_cast_5D882(0);
				_sv2v_jump = 2'b11;
			end
		end
	endfunction
	function automatic fpnew_pkg_is_first_enabled_multi;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:467:51
		input reg [2:0] fmt;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:468:51
		input reg [9:0] types;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:469:51
		input reg [0:4] cfg;
		reg [0:1] _sv2v_jump;
		begin
			_sv2v_jump = 2'b00;
			// Trace: core/cvfpu/src/fpnew_pkg.sv:470:5
			begin : sv2v_autoblock_7
				// Trace: core/cvfpu/src/fpnew_pkg.sv:470:10
				reg [31:0] i;
				// Trace: core/cvfpu/src/fpnew_pkg.sv:470:10
				begin : sv2v_autoblock_8
					reg [31:0] _sv2v_value_on_break;
					for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
						if (_sv2v_jump < 2'b10) begin
							_sv2v_jump = 2'b00;
							// Trace: core/cvfpu/src/fpnew_pkg.sv:471:7
							if (cfg[i] && (types[(4 - i) * 2+:2] == 2'd2)) begin
								fpnew_pkg_is_first_enabled_multi = sv2v_cast_5D882(i) == fmt;
								_sv2v_jump = 2'b11;
							end
							_sv2v_value_on_break = i;
						end
					if (!(_sv2v_jump < 2'b10))
						i = _sv2v_value_on_break;
					if (_sv2v_jump != 2'b11)
						_sv2v_jump = 2'b00;
				end
			end
			if (_sv2v_jump == 2'b00) begin
				fpnew_pkg_is_first_enabled_multi = 1'b0;
				_sv2v_jump = 2'b11;
			end
		end
	endfunction
	function automatic [31:0] fpnew_pkg_num_lanes;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:390:45
		input reg [31:0] width;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:390:65
		input reg [2:0] fmt;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:390:82
		input reg vec;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:391:5
		fpnew_pkg_num_lanes = (vec ? width / fpnew_pkg_fp_width(fmt) : 1);
	endfunction
	function automatic signed [31:0] sv2v_cast_32_signed;
		input reg signed [31:0] inp;
		sv2v_cast_32_signed = inp;
	endfunction
	function automatic [TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1:0] sv2v_cast_7CA2E;
		input reg [TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1:0] inp;
		sv2v_cast_7CA2E = inp;
	endfunction
	generate
		for (_gv_fmt_9 = 0; _gv_fmt_9 < sv2v_cast_32_signed(NUM_FORMATS); _gv_fmt_9 = _gv_fmt_9 + 1) begin : gen_parallel_slices
			localparam fmt = _gv_fmt_9;
			// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:88:5
			localparam [0:0] ANY_MERGED = fpnew_pkg_any_enabled_multi(FmtUnitTypes, FpFmtMask);
			// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:89:5
			localparam [0:0] IS_FIRST_MERGED = fpnew_pkg_is_first_enabled_multi(sv2v_cast_5D882(fmt), FmtUnitTypes, FpFmtMask);
			if (FpFmtMask[fmt] && (FmtUnitTypes[(4 - fmt) * 2+:2] == 2'd1)) begin : active_format
				// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:95:7
				wire in_valid;
				// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:97:7
				assign in_valid = in_valid_i & (dst_fmt_i == fmt);
				// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:100:7
				localparam [31:0] INTERNAL_LANES = fpnew_pkg_num_lanes(Width, sv2v_cast_5D882(fmt), EnableVectors);
				// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:101:7
				reg [INTERNAL_LANES - 1:0] mask_slice;
				// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:102:7
				always @(*) begin : sv2v_autoblock_9
					// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:102:24
					reg signed [31:0] b;
					if (_sv2v_0)
						;
					// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:102:24
					for (b = 0; b < INTERNAL_LANES; b = b + 1)
						begin
							// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:102:60
							mask_slice[b] = simd_mask_i[(NUM_LANES / INTERNAL_LANES) * b];
						end
				end
				// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:104:7
				fpnew_opgroup_fmt_slice_B2D7F_8C3BC #(
					.TagType_TagType_TagType_CVA6Cfg(TagType_TagType_CVA6Cfg),
					.TagType_TagType_TagType_config_pkg_NrMaxRules(TagType_TagType_config_pkg_NrMaxRules),
					.OpGroup(OpGroup),
					.FpFormat(sv2v_cast_5D882(fmt)),
					.Width(Width),
					.EnableVectors(EnableVectors),
					.NumPipeRegs(FmtPipeRegs[(4 - fmt) * 32+:32]),
					.PipeConfig(PipeConfig),
					.TrueSIMDClass(TrueSIMDClass)
				) i_fmt_slice(
					.clk_i(clk_i),
					.rst_ni(rst_ni),
					.operands_i(operands_i),
					.is_boxed_i(is_boxed_i[fmt * NUM_OPERANDS+:NUM_OPERANDS]),
					.rnd_mode_i(rnd_mode_i),
					.op_i(op_i),
					.op_mod_i(op_mod_i),
					.vectorial_op_i(vectorial_op_i),
					.tag_i(tag_i),
					.simd_mask_i(mask_slice),
					.in_valid_i(in_valid),
					.in_ready_o(fmt_in_ready[fmt]),
					.flush_i(flush_i),
					.result_o(fmt_outputs[(fmt * ((Width + 6) + TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)])) + (Width + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 5))-:((Width + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 5)) >= (6 + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0)) ? ((Width + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 5)) - (6 + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0))) + 1 : ((6 + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0)) - (Width + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 5))) + 1)]),
					.status_o(fmt_outputs[(fmt * ((Width + 6) + TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)])) + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 5)-:((TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 5) >= (1 + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0)) ? ((TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 5) - (1 + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0))) + 1 : ((1 + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0)) - (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 5)) + 1)]),
					.extension_bit_o(fmt_outputs[(fmt * ((Width + 6) + TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)])) + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0)]),
					.tag_o(fmt_outputs[(fmt * ((Width + 6) + TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)])) + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1)-:TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]]),
					.out_valid_o(fmt_out_valid[fmt]),
					.out_ready_i(fmt_out_ready[fmt]),
					.busy_o(fmt_busy[fmt])
				);
			end
			else if ((FpFmtMask[fmt] && ANY_MERGED) && !IS_FIRST_MERGED) begin : merged_unused
				// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:138:7
				localparam FMT = fpnew_pkg_get_first_enabled_multi(FmtUnitTypes, FpFmtMask);
				// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:140:7
				assign fmt_in_ready[fmt] = fmt_in_ready[sv2v_cast_32_signed(FMT)];
				// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:142:7
				assign fmt_out_valid[fmt] = 1'b0;
				// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:143:7
				assign fmt_busy[fmt] = 1'b0;
				// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:145:7
				assign fmt_outputs[(fmt * ((Width + 6) + TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)])) + (Width + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 5))-:((Width + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 5)) >= (6 + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0)) ? ((Width + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 5)) - (6 + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0))) + 1 : ((6 + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0)) - (Width + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 5))) + 1)] = {Width {fpnew_pkg_DONT_CARE}};
				// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:146:7
				assign fmt_outputs[(fmt * ((Width + 6) + TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)])) + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 5)-:((TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 5) >= (1 + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0)) ? ((TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 5) - (1 + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0))) + 1 : ((1 + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0)) - (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 5)) + 1)] = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
				// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:147:7
				assign fmt_outputs[(fmt * ((Width + 6) + TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)])) + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0)] = fpnew_pkg_DONT_CARE;
				// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:148:7
				assign fmt_outputs[(fmt * ((Width + 6) + TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)])) + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1)-:TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]] = sv2v_cast_7CA2E(fpnew_pkg_DONT_CARE);
			end
			else if (!FpFmtMask[fmt] || (FmtUnitTypes[(4 - fmt) * 2+:2] == 2'd0)) begin : disable_fmt
				// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:152:7
				assign fmt_in_ready[fmt] = 1'b0;
				// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:153:7
				assign fmt_out_valid[fmt] = 1'b0;
				// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:154:7
				assign fmt_busy[fmt] = 1'b0;
				// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:156:7
				assign fmt_outputs[(fmt * ((Width + 6) + TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)])) + (Width + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 5))-:((Width + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 5)) >= (6 + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0)) ? ((Width + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 5)) - (6 + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0))) + 1 : ((6 + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0)) - (Width + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 5))) + 1)] = {Width {fpnew_pkg_DONT_CARE}};
				// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:157:7
				assign fmt_outputs[(fmt * ((Width + 6) + TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)])) + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 5)-:((TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 5) >= (1 + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0)) ? ((TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 5) - (1 + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0))) + 1 : ((1 + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0)) - (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 5)) + 1)] = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
				// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:158:7
				assign fmt_outputs[(fmt * ((Width + 6) + TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)])) + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0)] = fpnew_pkg_DONT_CARE;
				// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:159:7
				assign fmt_outputs[(fmt * ((Width + 6) + TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)])) + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1)-:TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]] = sv2v_cast_7CA2E(fpnew_pkg_DONT_CARE);
			end
		end
	endgenerate
	// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:166:3
	function automatic [31:0] fpnew_pkg_get_num_regs_multi;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:485:54
		input reg [159:0] regs;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:486:54
		input reg [9:0] types;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:487:54
		input reg [0:4] cfg;
		// Trace: core/cvfpu/src/fpnew_pkg.sv:488:5
		reg [31:0] res;
		begin
			res = 0;
			// Trace: core/cvfpu/src/fpnew_pkg.sv:489:5
			begin : sv2v_autoblock_10
				// Trace: core/cvfpu/src/fpnew_pkg.sv:489:10
				reg [31:0] i;
				// Trace: core/cvfpu/src/fpnew_pkg.sv:489:10
				for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
					begin
						// Trace: core/cvfpu/src/fpnew_pkg.sv:490:7
						if (cfg[i] && (types[(4 - i) * 2+:2] == 2'd2))
							// Trace: core/cvfpu/src/fpnew_pkg.sv:490:41
							res = fpnew_pkg_maximum(res, regs[(4 - i) * 32+:32]);
					end
			end
			fpnew_pkg_get_num_regs_multi = res;
		end
	endfunction
	generate
		if (fpnew_pkg_any_enabled_multi(FmtUnitTypes, FpFmtMask)) begin : gen_merged_slice
			// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:168:5
			localparam FMT = fpnew_pkg_get_first_enabled_multi(FmtUnitTypes, FpFmtMask);
			// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:169:5
			localparam REG = fpnew_pkg_get_num_regs_multi(FmtPipeRegs, FmtUnitTypes, FpFmtMask);
			// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:171:5
			wire in_valid;
			// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:173:5
			assign in_valid = in_valid_i & (FmtUnitTypes[(4 - dst_fmt_i) * 2+:2] == 2'd2);
			// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:175:5
			fpnew_opgroup_multifmt_slice_983D9_76A82 #(
				.TagType_TagType_TagType_CVA6Cfg(TagType_TagType_CVA6Cfg),
				.TagType_TagType_TagType_config_pkg_NrMaxRules(TagType_TagType_config_pkg_NrMaxRules),
				.OpGroup(OpGroup),
				.Width(Width),
				.FpFmtConfig(FpFmtMask),
				.IntFmtConfig(IntFmtMask),
				.EnableVectors(EnableVectors),
				.NumPipeRegs(REG),
				.PipeConfig(PipeConfig)
			) i_multifmt_slice(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.operands_i(operands_i),
				.is_boxed_i(is_boxed_i),
				.rnd_mode_i(rnd_mode_i),
				.op_i(op_i),
				.op_mod_i(op_mod_i),
				.src_fmt_i(src_fmt_i),
				.dst_fmt_i(dst_fmt_i),
				.int_fmt_i(int_fmt_i),
				.vectorial_op_i(vectorial_op_i),
				.tag_i(tag_i),
				.simd_mask_i(simd_mask_i),
				.in_valid_i(in_valid),
				.in_ready_o(fmt_in_ready[FMT]),
				.flush_i(flush_i),
				.result_o(fmt_outputs[(FMT * ((Width + 6) + TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)])) + (Width + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 5))-:((Width + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 5)) >= (6 + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0)) ? ((Width + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 5)) - (6 + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0))) + 1 : ((6 + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0)) - (Width + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 5))) + 1)]),
				.status_o(fmt_outputs[(FMT * ((Width + 6) + TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)])) + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 5)-:((TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 5) >= (1 + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0)) ? ((TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 5) - (1 + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0))) + 1 : ((1 + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0)) - (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 5)) + 1)]),
				.extension_bit_o(fmt_outputs[(FMT * ((Width + 6) + TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)])) + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0)]),
				.tag_o(fmt_outputs[(FMT * ((Width + 6) + TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)])) + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1)-:TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]]),
				.out_valid_o(fmt_out_valid[FMT]),
				.out_ready_i(fmt_out_ready[FMT]),
				.busy_o(fmt_busy[FMT])
			);
		end
	endgenerate
	// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:215:3
	wire [((Width + 6) + TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) - 1:0] arbiter_output;
	// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:218:3
	localparam [31:0] sv2v_uu_i_arbiter_NumIn = NUM_FORMATS;
	localparam [31:0] sv2v_uu_i_arbiter_IdxWidth = $unsigned(3);
	// removed localparam type sv2v_uu_i_arbiter_rr_i
	localparam [sv2v_uu_i_arbiter_IdxWidth - 1:0] sv2v_uu_i_arbiter_ext_rr_i_0 = 1'sb0;
	rr_arb_tree_11E95_B691C #(
		.DataType_TagType_TagType_CVA6Cfg(TagType_TagType_CVA6Cfg),
		.DataType_TagType_TagType_config_pkg_NrMaxRules(TagType_TagType_config_pkg_NrMaxRules),
		.DataType_Width(Width),
		.NumIn(NUM_FORMATS),
		.AxiVldRdy(1'b1)
	) i_arbiter(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(flush_i),
		.rr_i(sv2v_uu_i_arbiter_ext_rr_i_0),
		.req_i(fmt_out_valid),
		.gnt_o(fmt_out_ready),
		.data_i(fmt_outputs),
		.gnt_i(out_ready_i),
		.req_o(out_valid_o),
		.data_o(arbiter_output),
		.idx_o()
	);
	// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:237:3
	assign result_o = arbiter_output[Width + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 5)-:((Width + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 5)) >= (6 + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0)) ? ((Width + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 5)) - (6 + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0))) + 1 : ((6 + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0)) - (Width + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 5))) + 1)];
	// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:238:3
	assign status_o = arbiter_output[TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 5-:((TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 5) >= (1 + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0)) ? ((TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 5) - (1 + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0))) + 1 : ((1 + (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0)) - (TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 5)) + 1)];
	// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:239:3
	assign extension_bit_o = arbiter_output[TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0];
	// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:240:3
	assign tag_o = arbiter_output[TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1-:TagType_TagType_CVA6Cfg[8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))-:((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353))))))))) - (8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((8910 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1354))))))))) - (8942 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + (32 + ((TagType_TagType_config_pkg_NrMaxRules * 64) + ((TagType_TagType_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]];
	// Trace: core/cvfpu/src/fpnew_opgroup_block.sv:242:3
	assign busy_o = |fmt_busy;
	initial _sv2v_0 = 0;
endmodule
