module btb_C3780_5CA66 (
	clk_i,
	rst_ni,
	flush_bp_i,
	debug_mode_i,
	vpc_i,
	btb_update_i,
	btb_prediction_o
);
	// removed localparam type btb_prediction_t_CVA6Cfg_type
	// removed localparam type btb_prediction_t_config_pkg_NrMaxRules_type
	parameter [17102:0] btb_prediction_t_CVA6Cfg = 0;
	parameter signed [31:0] btb_prediction_t_config_pkg_NrMaxRules = 0;
	// removed localparam type btb_update_t_CVA6Cfg_type
	// removed localparam type btb_update_t_config_pkg_NrMaxRules_type
	parameter [17102:0] btb_update_t_CVA6Cfg = 0;
	parameter signed [31:0] btb_update_t_config_pkg_NrMaxRules = 0;
	reg _sv2v_0;
	// Trace: core/frontend/btb.sv:29:15
	localparam config_pkg_NrMaxRules = 16;
	// removed localparam type config_pkg_cache_type_t
	// removed localparam type config_pkg_noc_type_e
	// removed localparam type config_pkg_vm_mode_t
	// removed localparam type config_pkg_cva6_cfg_t
	localparam [17102:0] config_pkg_cva6_cfg_empty = 17103'd0;
	parameter [17102:0] CVA6Cfg = config_pkg_cva6_cfg_empty;
	// Trace: core/frontend/btb.sv:30:20
	// removed localparam type btb_update_t
	// Trace: core/frontend/btb.sv:31:20
	// removed localparam type btb_prediction_t
	// Trace: core/frontend/btb.sv:32:15
	parameter signed [31:0] NR_ENTRIES = 8;
	// Trace: core/frontend/btb.sv:35:5
	input wire clk_i;
	// Trace: core/frontend/btb.sv:37:5
	input wire rst_ni;
	// Trace: core/frontend/btb.sv:39:5
	input wire flush_bp_i;
	// Trace: core/frontend/btb.sv:41:5
	input wire debug_mode_i;
	// Trace: core/frontend/btb.sv:43:5
	input wire [CVA6Cfg[17070-:32] - 1:0] vpc_i;
	// Trace: core/frontend/btb.sv:45:5
	input wire [((1 + btb_update_t_CVA6Cfg[9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + btb_update_t_CVA6Cfg[9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) - 1:0] btb_update_i;
	// Trace: core/frontend/btb.sv:47:5
	output wire [(CVA6Cfg[579-:32] * (1 + btb_prediction_t_CVA6Cfg[9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)])) - 1:0] btb_prediction_o;
	// Trace: core/frontend/btb.sv:50:3
	localparam OFFSET = (CVA6Cfg[16544] == 1'b1 ? 1 : 2);
	// Trace: core/frontend/btb.sv:52:3
	localparam NR_ROWS = NR_ENTRIES / CVA6Cfg[579-:32];
	// Trace: core/frontend/btb.sv:54:3
	localparam ROW_ADDR_BITS = $clog2(CVA6Cfg[579-:32]);
	// Trace: core/frontend/btb.sv:55:3
	localparam ROW_INDEX_BITS = (CVA6Cfg[16544] == 1'b1 ? $clog2(CVA6Cfg[579-:32]) : 1);
	// Trace: core/frontend/btb.sv:57:3
	localparam PREDICTION_BITS = ($clog2(NR_ROWS) + OFFSET) + ROW_ADDR_BITS;
	// Trace: core/frontend/btb.sv:59:3
	localparam ANTIALIAS_BITS = 8;
	// Trace: core/frontend/btb.sv:61:3
	localparam BRAM_WORD_BITS = 1 + btb_prediction_t_CVA6Cfg[9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)];
	// Trace: core/frontend/btb.sv:63:3
	unread i_unread(.d_i(|vpc_i));
	// Trace: core/frontend/btb.sv:66:3
	wire [$clog2(NR_ROWS) - 1:0] index;
	wire [$clog2(NR_ROWS) - 1:0] update_pc;
	// Trace: core/frontend/btb.sv:67:3
	wire [ROW_INDEX_BITS - 1:0] update_row_index;
	// Trace: core/frontend/btb.sv:69:3
	assign index = vpc_i[PREDICTION_BITS - 1:ROW_ADDR_BITS + OFFSET];
	// Trace: core/frontend/btb.sv:70:3
	assign update_pc = btb_update_i[(btb_update_t_CVA6Cfg[9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (btb_update_t_CVA6Cfg[9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1)) - ((btb_update_t_CVA6Cfg[9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1) - (PREDICTION_BITS - 1)):(btb_update_t_CVA6Cfg[9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (btb_update_t_CVA6Cfg[9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1)) - ((btb_update_t_CVA6Cfg[9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1) - (ROW_ADDR_BITS + OFFSET))];
	// Trace: core/frontend/btb.sv:71:3
	generate
		if (CVA6Cfg[16544]) begin : gen_update_row_index
			// Trace: core/frontend/btb.sv:72:5
			assign update_row_index = btb_update_i[(btb_update_t_CVA6Cfg[9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (btb_update_t_CVA6Cfg[9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1)) - ((btb_update_t_CVA6Cfg[9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1) - ((ROW_ADDR_BITS + OFFSET) - 1)):(btb_update_t_CVA6Cfg[9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (btb_update_t_CVA6Cfg[9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1)) - ((btb_update_t_CVA6Cfg[9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1) - OFFSET)];
		end
		else begin : genblk1
			// Trace: core/frontend/btb.sv:74:5
			assign update_row_index = 1'sb0;
		end
	endgenerate
	// Trace: core/frontend/btb.sv:77:3
	function automatic [(1 + btb_prediction_t_CVA6Cfg[9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) - 1:0] sv2v_cast_ABDD7;
		input reg [(1 + btb_prediction_t_CVA6Cfg[9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) - 1:0] inp;
		sv2v_cast_ABDD7 = inp;
	endfunction
	generate
		if (CVA6Cfg[16876]) begin : gen_fpga_btb
			// Trace: core/frontend/btb.sv:78:5
			wire [CVA6Cfg[579-:32] - 1:0] btb_ram_csel_prediction;
			// Trace: core/frontend/btb.sv:79:5
			wire [CVA6Cfg[579-:32] - 1:0] btb_ram_we_prediction;
			// Trace: core/frontend/btb.sv:80:5
			wire [(CVA6Cfg[579-:32] * $clog2(NR_ROWS)) - 1:0] btb_ram_addr_prediction;
			// Trace: core/frontend/btb.sv:81:5
			wire [(CVA6Cfg[579-:32] * BRAM_WORD_BITS) - 1:0] btb_ram_wdata_prediction;
			// Trace: core/frontend/btb.sv:82:5
			wire [(CVA6Cfg[579-:32] * BRAM_WORD_BITS) - 1:0] btb_ram_rdata_prediction;
			// Trace: core/frontend/btb.sv:84:5
			reg [CVA6Cfg[579-:32] - 1:0] btb_ram_csel_update;
			// Trace: core/frontend/btb.sv:85:5
			reg [CVA6Cfg[579-:32] - 1:0] btb_ram_we_update;
			// Trace: core/frontend/btb.sv:86:5
			reg [(CVA6Cfg[579-:32] * $clog2(NR_ROWS)) - 1:0] btb_ram_addr_update;
			// Trace: core/frontend/btb.sv:87:5
			reg [(CVA6Cfg[579-:32] * BRAM_WORD_BITS) - 1:0] btb_ram_wdata_update;
			genvar _gv_i_54;
			for (_gv_i_54 = 0; _gv_i_54 < CVA6Cfg[579-:32]; _gv_i_54 = _gv_i_54 + 1) begin : gen_btb_output
				localparam i = _gv_i_54;
				// Trace: core/frontend/btb.sv:91:7
				assign btb_ram_csel_prediction[i] = 1'b1;
				// Trace: core/frontend/btb.sv:92:7
				assign btb_ram_we_prediction[i] = 1'b0;
				// Trace: core/frontend/btb.sv:93:7
				assign btb_ram_wdata_prediction = 1'sb0;
				// Trace: core/frontend/btb.sv:94:7
				assign btb_ram_addr_prediction[i * $clog2(NR_ROWS)+:$clog2(NR_ROWS)] = index;
				// Trace: core/frontend/btb.sv:95:7
				assign btb_prediction_o[i * (1 + btb_prediction_t_CVA6Cfg[9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)])+:1 + btb_prediction_t_CVA6Cfg[9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]] = btb_ram_rdata_prediction[i * BRAM_WORD_BITS+:BRAM_WORD_BITS];
			end
			// Trace: core/frontend/btb.sv:102:5
			always @(*) begin : update_branch_predict
				if (_sv2v_0)
					;
				// Trace: core/frontend/btb.sv:103:7
				btb_ram_csel_update = 1'sb0;
				// Trace: core/frontend/btb.sv:104:7
				btb_ram_we_update = 1'sb0;
				// Trace: core/frontend/btb.sv:105:7
				btb_ram_addr_update = 1'sb0;
				// Trace: core/frontend/btb.sv:106:7
				btb_ram_wdata_update = 1'sb0;
				// Trace: core/frontend/btb.sv:108:7
				if (btb_update_i[1 + (btb_update_t_CVA6Cfg[9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (btb_update_t_CVA6Cfg[9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1))] && !debug_mode_i)
					// Trace: core/frontend/btb.sv:109:9
					begin : sv2v_autoblock_1
						// Trace: core/frontend/btb.sv:109:14
						reg signed [31:0] i;
						// Trace: core/frontend/btb.sv:109:14
						for (i = 0; i < CVA6Cfg[579-:32]; i = i + 1)
							begin
								// Trace: core/frontend/btb.sv:110:11
								if (update_row_index == i) begin
									// Trace: core/frontend/btb.sv:111:13
									btb_ram_csel_update[i] = 1'b1;
									// Trace: core/frontend/btb.sv:112:13
									btb_ram_we_update[i] = 1'b1;
									// Trace: core/frontend/btb.sv:113:13
									btb_ram_addr_update[i * $clog2(NR_ROWS)+:$clog2(NR_ROWS)] = update_pc;
									// Trace: core/frontend/btb.sv:114:13
									btb_ram_wdata_update[i * BRAM_WORD_BITS+:BRAM_WORD_BITS] = {1'b1, btb_update_i[btb_update_t_CVA6Cfg[9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1-:btb_update_t_CVA6Cfg[9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]]};
								end
							end
					end
			end
			genvar _gv_i_55;
			for (_gv_i_55 = 0; _gv_i_55 < CVA6Cfg[579-:32]; _gv_i_55 = _gv_i_55 + 1) begin : gen_btb_ram
				localparam i = _gv_i_55;
				// Trace: core/frontend/btb.sv:123:7
				SyncDpRam #(
					.ADDR_WIDTH($clog2(NR_ROWS)),
					.DATA_DEPTH(NR_ROWS),
					.DATA_WIDTH(BRAM_WORD_BITS),
					.OUT_REGS(0),
					.SIM_INIT(1)
				) i_btb_ram(
					.Clk_CI(clk_i),
					.Rst_RBI(rst_ni),
					.CSelA_SI(btb_ram_csel_update[i]),
					.WrEnA_SI(btb_ram_we_update[i]),
					.AddrA_DI(btb_ram_addr_update[i * $clog2(NR_ROWS)+:$clog2(NR_ROWS)]),
					.WrDataA_DI(btb_ram_wdata_update[i * BRAM_WORD_BITS+:BRAM_WORD_BITS]),
					.RdDataA_DO(),
					.CSelB_SI(btb_ram_csel_prediction[i]),
					.WrEnB_SI(btb_ram_we_prediction[i]),
					.AddrB_DI(btb_ram_addr_prediction[i * $clog2(NR_ROWS)+:$clog2(NR_ROWS)]),
					.WrDataB_DI(btb_ram_wdata_prediction[i * BRAM_WORD_BITS+:BRAM_WORD_BITS]),
					.RdDataB_DO(btb_ram_rdata_prediction[i * BRAM_WORD_BITS+:BRAM_WORD_BITS])
				);
			end
		end
		else begin : gen_asic_btb
			// Trace: core/frontend/btb.sv:151:5
			reg [((NR_ROWS * CVA6Cfg[579-:32]) * (1 + btb_prediction_t_CVA6Cfg[9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)])) - 1:0] btb_d;
			reg [((NR_ROWS * CVA6Cfg[579-:32]) * (1 + btb_prediction_t_CVA6Cfg[9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)])) - 1:0] btb_q;
			genvar _gv_i_56;
			for (_gv_i_56 = 0; _gv_i_56 < CVA6Cfg[579-:32]; _gv_i_56 = _gv_i_56 + 1) begin : gen_btb_output
				localparam i = _gv_i_56;
				// Trace: core/frontend/btb.sv:157:7
				assign btb_prediction_o[i * (1 + btb_prediction_t_CVA6Cfg[9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)])+:1 + btb_prediction_t_CVA6Cfg[9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]] = btb_q[((index * CVA6Cfg[579-:32]) + i) * (1 + btb_prediction_t_CVA6Cfg[9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)])+:1 + btb_prediction_t_CVA6Cfg[9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]];
			end
			// Trace: core/frontend/btb.sv:164:5
			always @(*) begin : update_branch_predict
				if (_sv2v_0)
					;
				// Trace: core/frontend/btb.sv:165:7
				btb_d = btb_q;
				// Trace: core/frontend/btb.sv:167:7
				if (btb_update_i[1 + (btb_update_t_CVA6Cfg[9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (btb_update_t_CVA6Cfg[9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1))] && !debug_mode_i) begin
					// Trace: core/frontend/btb.sv:168:9
					btb_d[(((update_pc * CVA6Cfg[579-:32]) + update_row_index) * (1 + btb_prediction_t_CVA6Cfg[9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)])) + (btb_prediction_t_CVA6Cfg[9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0)] = 1'b1;
					// Trace: core/frontend/btb.sv:170:9
					btb_d[(((update_pc * CVA6Cfg[579-:32]) + update_row_index) * (1 + btb_prediction_t_CVA6Cfg[9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)])) + (btb_prediction_t_CVA6Cfg[9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1)-:btb_prediction_t_CVA6Cfg[9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]] = btb_update_i[btb_update_t_CVA6Cfg[9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] - 1-:btb_update_t_CVA6Cfg[9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_update_t_config_pkg_NrMaxRules * 64) + ((btb_update_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]];
				end
			end
			// Trace: core/frontend/btb.sv:175:5
			always @(posedge clk_i or negedge rst_ni)
				// Trace: core/frontend/btb.sv:176:7
				if (!rst_ni)
					// Trace: core/frontend/btb.sv:178:9
					begin : sv2v_autoblock_2
						// Trace: core/frontend/btb.sv:178:14
						reg signed [31:0] i;
						// Trace: core/frontend/btb.sv:178:14
						for (i = 0; i < NR_ROWS; i = i + 1)
							begin
								// Trace: core/frontend/btb.sv:178:43
								btb_q[(1 + btb_prediction_t_CVA6Cfg[9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) * (i * CVA6Cfg[579-:32])+:(1 + btb_prediction_t_CVA6Cfg[9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) * CVA6Cfg[579-:32]] <= {CVA6Cfg[579-:32] {sv2v_cast_ABDD7(0)}};
							end
					end
				else
					// Trace: core/frontend/btb.sv:181:9
					if (flush_bp_i)
						// Trace: core/frontend/btb.sv:182:11
						begin : sv2v_autoblock_3
							// Trace: core/frontend/btb.sv:182:16
							reg signed [31:0] i;
							// Trace: core/frontend/btb.sv:182:16
							for (i = 0; i < NR_ROWS; i = i + 1)
								begin
									// Trace: core/frontend/btb.sv:183:13
									begin : sv2v_autoblock_4
										// Trace: core/frontend/btb.sv:183:18
										reg signed [31:0] j;
										// Trace: core/frontend/btb.sv:183:18
										for (j = 0; j < CVA6Cfg[579-:32]; j = j + 1)
											begin
												// Trace: core/frontend/btb.sv:184:15
												btb_q[(((i * CVA6Cfg[579-:32]) + j) * (1 + btb_prediction_t_CVA6Cfg[9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)])) + (btb_prediction_t_CVA6Cfg[9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9477 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9509 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + (32 + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + ((btb_prediction_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0)] <= 1'b0;
											end
									end
								end
						end
					else
						// Trace: core/frontend/btb.sv:188:11
						btb_q <= btb_d;
		end
	endgenerate
	initial _sv2v_0 = 0;
endmodule
