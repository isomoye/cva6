module scoreboard_20CF9_053D6 (
	clk_i,
	rst_ni,
	sb_full_o,
	flush_unissued_instr_i,
	flush_i,
	rd_clobber_gpr_o,
	rd_clobber_fpr_o,
	x_transaction_accepted_i,
	x_issue_writeback_i,
	x_id_i,
	rs1_i,
	rs1_o,
	rs1_valid_o,
	rs2_i,
	rs2_o,
	rs2_valid_o,
	rs3_i,
	rs3_o,
	rs3_valid_o,
	commit_instr_o,
	commit_drop_o,
	commit_ack_i,
	decoded_instr_i,
	orig_instr_i,
	decoded_instr_valid_i,
	decoded_instr_ack_o,
	issue_instr_o,
	orig_instr_o,
	issue_instr_valid_o,
	issue_ack_i,
	resolved_branch_i,
	trans_id_i,
	wbdata_i,
	ex_i,
	wt_valid_i,
	x_we_i,
	x_rd_i,
	rvfi_issue_pointer_o,
	rvfi_commit_pointer_o
);
	// removed localparam type bp_resolve_t_bp_resolve_t_CVA6Cfg_type
	parameter [17102:0] bp_resolve_t_bp_resolve_t_CVA6Cfg = 0;
	// removed localparam type exception_t_exception_t_CVA6Cfg_type
	parameter [17102:0] exception_t_exception_t_CVA6Cfg = 0;
	// removed localparam type rs3_len_t_CVA6Cfg_type
	parameter [17102:0] rs3_len_t_CVA6Cfg = 0;
	// removed localparam type scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg_type
	parameter [17102:0] scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg = 0;
	reg _sv2v_0;
	// Trace: core/scoreboard.sv:16:15
	localparam config_pkg_NrMaxRules = 16;
	// removed localparam type config_pkg_cache_type_t
	// removed localparam type config_pkg_noc_type_e
	// removed localparam type config_pkg_vm_mode_t
	// removed localparam type config_pkg_cva6_cfg_t
	localparam [17102:0] config_pkg_cva6_cfg_empty = 17103'd0;
	parameter [17102:0] CVA6Cfg = config_pkg_cva6_cfg_empty;
	// Trace: core/scoreboard.sv:17:20
	// removed localparam type bp_resolve_t
	// Trace: core/scoreboard.sv:18:20
	// removed localparam type exception_t
	// Trace: core/scoreboard.sv:19:20
	// removed localparam type scoreboard_entry_t
	// Trace: core/scoreboard.sv:20:20
	// removed localparam type rs3_len_t
	// Trace: core/scoreboard.sv:23:5
	input wire clk_i;
	// Trace: core/scoreboard.sv:25:5
	input wire rst_ni;
	// Trace: core/scoreboard.sv:27:5
	output wire sb_full_o;
	// Trace: core/scoreboard.sv:29:5
	input wire flush_unissued_instr_i;
	// Trace: core/scoreboard.sv:31:5
	input wire flush_i;
	// Trace: core/scoreboard.sv:33:5
	localparam ariane_pkg_REG_ADDR_SIZE = 5;
	// removed localparam type ariane_pkg_fu_t
	output wire [127:0] rd_clobber_gpr_o;
	// Trace: core/scoreboard.sv:35:5
	output wire [127:0] rd_clobber_fpr_o;
	// Trace: core/scoreboard.sv:37:5
	input wire x_transaction_accepted_i;
	// Trace: core/scoreboard.sv:38:5
	input wire x_issue_writeback_i;
	// Trace: core/scoreboard.sv:39:5
	input wire [CVA6Cfg[16503-:32] - 1:0] x_id_i;
	// Trace: core/scoreboard.sv:41:5
	input wire [(CVA6Cfg[16841-:32] * 5) - 1:0] rs1_i;
	// Trace: core/scoreboard.sv:43:5
	output wire [(CVA6Cfg[16841-:32] * CVA6Cfg[17102-:32]) - 1:0] rs1_o;
	// Trace: core/scoreboard.sv:45:5
	output wire [CVA6Cfg[16841-:32] - 1:0] rs1_valid_o;
	// Trace: core/scoreboard.sv:48:5
	input wire [(CVA6Cfg[16841-:32] * 5) - 1:0] rs2_i;
	// Trace: core/scoreboard.sv:50:5
	output wire [(CVA6Cfg[16841-:32] * CVA6Cfg[17102-:32]) - 1:0] rs2_o;
	// Trace: core/scoreboard.sv:52:5
	output wire [CVA6Cfg[16841-:32] - 1:0] rs2_valid_o;
	// Trace: core/scoreboard.sv:55:5
	input wire [(CVA6Cfg[16841-:32] * 5) - 1:0] rs3_i;
	// Trace: core/scoreboard.sv:57:5
	output wire [(CVA6Cfg[16841-:32] * (rs3_len_t_CVA6Cfg[16433-:32] == 3 ? rs3_len_t_CVA6Cfg[17102-:32] : rs3_len_t_CVA6Cfg[16469-:32])) - 1:0] rs3_o;
	// Trace: core/scoreboard.sv:59:5
	output wire [CVA6Cfg[16841-:32] - 1:0] rs3_valid_o;
	// Trace: core/scoreboard.sv:63:5
	output reg [((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (CVA6Cfg[16873-:32] * (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5)) - 1 : (CVA6Cfg[16873-:32] * (1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 3)):((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 0 : ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)] commit_instr_o;
	// Trace: core/scoreboard.sv:65:5
	output reg [CVA6Cfg[16873-:32] - 1:0] commit_drop_o;
	// Trace: core/scoreboard.sv:67:5
	input wire [CVA6Cfg[16873-:32] - 1:0] commit_ack_i;
	// Trace: core/scoreboard.sv:72:5
	input wire [((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (CVA6Cfg[16841-:32] * (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5)) - 1 : (CVA6Cfg[16841-:32] * (1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 3)):((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 0 : ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)] decoded_instr_i;
	// Trace: core/scoreboard.sv:74:5
	input wire [(CVA6Cfg[16841-:32] * 32) - 1:0] orig_instr_i;
	// Trace: core/scoreboard.sv:76:5
	input wire [CVA6Cfg[16841-:32] - 1:0] decoded_instr_valid_i;
	// Trace: core/scoreboard.sv:78:5
	output reg [CVA6Cfg[16841-:32] - 1:0] decoded_instr_ack_o;
	// Trace: core/scoreboard.sv:82:5
	output reg [((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (CVA6Cfg[16841-:32] * (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5)) - 1 : (CVA6Cfg[16841-:32] * (1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 3)):((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 0 : ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)] issue_instr_o;
	// Trace: core/scoreboard.sv:84:5
	output reg [(CVA6Cfg[16841-:32] * 32) - 1:0] orig_instr_o;
	// Trace: core/scoreboard.sv:86:5
	output reg [CVA6Cfg[16841-:32] - 1:0] issue_instr_valid_o;
	// Trace: core/scoreboard.sv:88:5
	input wire [CVA6Cfg[16841-:32] - 1:0] issue_ack_i;
	// Trace: core/scoreboard.sv:91:5
	input wire [((1 + bp_resolve_t_bp_resolve_t_CVA6Cfg[17070-:32]) + bp_resolve_t_bp_resolve_t_CVA6Cfg[17070-:32]) + 4:0] resolved_branch_i;
	// Trace: core/scoreboard.sv:93:5
	input wire [(CVA6Cfg[16401-:32] * CVA6Cfg[16503-:32]) - 1:0] trans_id_i;
	// Trace: core/scoreboard.sv:95:5
	input wire [(CVA6Cfg[16401-:32] * CVA6Cfg[17102-:32]) - 1:0] wbdata_i;
	// Trace: core/scoreboard.sv:97:5
	input wire [((((exception_t_exception_t_CVA6Cfg[17102-:32] + exception_t_exception_t_CVA6Cfg[17102-:32]) + exception_t_exception_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? (CVA6Cfg[16401-:32] * (((exception_t_exception_t_CVA6Cfg[17102-:32] + exception_t_exception_t_CVA6Cfg[17102-:32]) + exception_t_exception_t_CVA6Cfg[17006-:32]) + 34)) - 1 : (CVA6Cfg[16401-:32] * (1 - (((exception_t_exception_t_CVA6Cfg[17102-:32] + exception_t_exception_t_CVA6Cfg[17102-:32]) + exception_t_exception_t_CVA6Cfg[17006-:32]) + 33))) + (((exception_t_exception_t_CVA6Cfg[17102-:32] + exception_t_exception_t_CVA6Cfg[17102-:32]) + exception_t_exception_t_CVA6Cfg[17006-:32]) + 32)):((((exception_t_exception_t_CVA6Cfg[17102-:32] + exception_t_exception_t_CVA6Cfg[17102-:32]) + exception_t_exception_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? 0 : ((exception_t_exception_t_CVA6Cfg[17102-:32] + exception_t_exception_t_CVA6Cfg[17102-:32]) + exception_t_exception_t_CVA6Cfg[17006-:32]) + 33)] ex_i;
	// Trace: core/scoreboard.sv:99:5
	input wire [CVA6Cfg[16401-:32] - 1:0] wt_valid_i;
	// Trace: core/scoreboard.sv:101:5
	input wire x_we_i;
	// Trace: core/scoreboard.sv:103:5
	input wire [4:0] x_rd_i;
	// Trace: core/scoreboard.sv:106:5
	output wire [(CVA6Cfg[16841-:32] * CVA6Cfg[16503-:32]) - 1:0] rvfi_issue_pointer_o;
	// Trace: core/scoreboard.sv:108:5
	output wire [(CVA6Cfg[16873-:32] * CVA6Cfg[16503-:32]) - 1:0] rvfi_commit_pointer_o;
	// Trace: core/scoreboard.sv:112:3
	// removed localparam type sb_mem_t
	// Trace: core/scoreboard.sv:118:3
	reg [(CVA6Cfg[16535-:32] * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) - 1:0] mem_q;
	reg [(CVA6Cfg[16535-:32] * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) - 1:0] mem_n;
	// Trace: core/scoreboard.sv:119:3
	wire [CVA6Cfg[16535-:32] - 1:0] still_issued;
	// Trace: core/scoreboard.sv:121:3
	wire [CVA6Cfg[16841-:32] - 1:0] issue_full;
	// Trace: core/scoreboard.sv:122:3
	wire [(2 * (CVA6Cfg[16535-:32] / 2)) - 1:0] issued_instrs_even_odd;
	// Trace: core/scoreboard.sv:124:3
	wire bmiss;
	// Trace: core/scoreboard.sv:125:3
	wire [CVA6Cfg[16503-:32] - 1:0] after_flu_wb;
	// Trace: core/scoreboard.sv:126:3
	wire [CVA6Cfg[16535-:32] - 1:0] speculative_instrs;
	// Trace: core/scoreboard.sv:128:3
	reg [CVA6Cfg[16841-:32] - 1:0] num_issue;
	// Trace: core/scoreboard.sv:129:3
	reg [CVA6Cfg[16503-:32] - 1:0] issue_pointer_n;
	reg [CVA6Cfg[16503-:32] - 1:0] issue_pointer_q;
	// Trace: core/scoreboard.sv:130:3
	wire [(CVA6Cfg[16841-:32] >= 0 ? ((CVA6Cfg[16841-:32] + 1) * CVA6Cfg[16503-:32]) - 1 : ((1 - CVA6Cfg[16841-:32]) * CVA6Cfg[16503-:32]) + ((CVA6Cfg[16841-:32] * CVA6Cfg[16503-:32]) - 1)):(CVA6Cfg[16841-:32] >= 0 ? 0 : CVA6Cfg[16841-:32] * CVA6Cfg[16503-:32])] issue_pointer;
	// Trace: core/scoreboard.sv:132:3
	wire [(CVA6Cfg[16873-:32] * CVA6Cfg[16503-:32]) - 1:0] commit_pointer_n;
	reg [(CVA6Cfg[16873-:32] * CVA6Cfg[16503-:32]) - 1:0] commit_pointer_q;
	// Trace: core/scoreboard.sv:133:3
	wire [$clog2(CVA6Cfg[16873-:32]):0] num_commit;
	// Trace: core/scoreboard.sv:135:3
	genvar _gv_i_47;
	generate
		for (_gv_i_47 = 0; _gv_i_47 < CVA6Cfg[16535-:32]; _gv_i_47 = _gv_i_47 + 1) begin : genblk1
			localparam i = _gv_i_47;
			// Trace: core/scoreboard.sv:136:5
			assign still_issued[i] = mem_q[(i * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + (2 + (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 0))] & ~mem_q[(i * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 1)];
		end
	endgenerate
	// Trace: core/scoreboard.sv:139:3
	genvar _gv_i_48;
	generate
		for (_gv_i_48 = 0; _gv_i_48 < CVA6Cfg[16535-:32]; _gv_i_48 = _gv_i_48 + 1) begin : genblk2
			localparam i = _gv_i_48;
			// Trace: core/scoreboard.sv:140:5
			assign issued_instrs_even_odd[((i % 2) * (CVA6Cfg[16535-:32] / 2)) + (i / 2)] = mem_q[(i * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + (2 + (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 0))];
		end
	endgenerate
	// Trace: core/scoreboard.sv:144:3
	assign issue_full[0] = &issued_instrs_even_odd[0+:CVA6Cfg[16535-:32] / 2] && &issued_instrs_even_odd[CVA6Cfg[16535-:32] / 2+:CVA6Cfg[16535-:32] / 2];
	// Trace: core/scoreboard.sv:145:3
	generate
		if (CVA6Cfg[16874]) begin : assign_issue_full
			// Trace: core/scoreboard.sv:148:5
			assign issue_full[1] = &issued_instrs_even_odd[0+:CVA6Cfg[16535-:32] / 2] || &issued_instrs_even_odd[CVA6Cfg[16535-:32] / 2+:CVA6Cfg[16535-:32] / 2];
		end
	endgenerate
	// Trace: core/scoreboard.sv:151:3
	assign sb_full_o = issue_full[0];
	// Trace: core/scoreboard.sv:154:3
	always @(*) begin : commit_ports
		if (_sv2v_0)
			;
		// Trace: core/scoreboard.sv:155:5
		begin : sv2v_autoblock_1
			// Trace: core/scoreboard.sv:155:10
			reg [31:0] i;
			// Trace: core/scoreboard.sv:155:10
			for (i = 0; i < CVA6Cfg[16873-:32]; i = i + 1)
				begin
					// Trace: core/scoreboard.sv:156:7
					commit_instr_o[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 0 : ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) + (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))+:((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))] = mem_q[(commit_pointer_q[i * CVA6Cfg[16503-:32]+:CVA6Cfg[16503-:32]] * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) - 1)-:((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))];
					// Trace: core/scoreboard.sv:157:7
					commit_instr_o[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))))) + ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) >= (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + 1)) - 1)-:((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) >= (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + 1)] = commit_pointer_q[i * CVA6Cfg[16503-:32]+:CVA6Cfg[16503-:32]];
					// Trace: core/scoreboard.sv:158:7
					commit_drop_o[i] = mem_q[(commit_pointer_q[i * CVA6Cfg[16503-:32]+:CVA6Cfg[16503-:32]] * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 1)];
				end
		end
	end
	// Trace: core/scoreboard.sv:162:3
	assign issue_pointer[(CVA6Cfg[16841-:32] >= 0 ? 0 : CVA6Cfg[16841-:32]) * CVA6Cfg[16503-:32]+:CVA6Cfg[16503-:32]] = issue_pointer_q;
	// Trace: core/scoreboard.sv:163:3
	genvar _gv_i_49;
	generate
		for (_gv_i_49 = 0; _gv_i_49 < CVA6Cfg[16841-:32]; _gv_i_49 = _gv_i_49 + 1) begin : genblk4
			localparam i = _gv_i_49;
			// Trace: core/scoreboard.sv:164:5
			assign issue_pointer[(CVA6Cfg[16841-:32] >= 0 ? i + 1 : CVA6Cfg[16841-:32] - (i + 1)) * CVA6Cfg[16503-:32]+:CVA6Cfg[16503-:32]] = issue_pointer[(CVA6Cfg[16841-:32] >= 0 ? i : CVA6Cfg[16841-:32] - i) * CVA6Cfg[16503-:32]+:CVA6Cfg[16503-:32]] + 'd1;
		end
	endgenerate
	// Trace: core/scoreboard.sv:168:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: core/scoreboard.sv:169:5
		issue_instr_o = decoded_instr_i;
		// Trace: core/scoreboard.sv:170:5
		orig_instr_o = orig_instr_i;
		// Trace: core/scoreboard.sv:171:5
		begin : sv2v_autoblock_2
			// Trace: core/scoreboard.sv:171:10
			reg [31:0] i;
			// Trace: core/scoreboard.sv:171:10
			for (i = 0; i < CVA6Cfg[16841-:32]; i = i + 1)
				begin
					// Trace: core/scoreboard.sv:173:7
					issue_instr_o[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))))) + ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) >= (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + 1)) - 1)-:((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) >= (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + 1)] = issue_pointer[(CVA6Cfg[16841-:32] >= 0 ? i : CVA6Cfg[16841-:32] - i) * CVA6Cfg[16503-:32]+:CVA6Cfg[16503-:32]];
					// Trace: core/scoreboard.sv:175:7
					issue_instr_valid_o[i] = decoded_instr_valid_i[i] & ~issue_full[i];
					// Trace: core/scoreboard.sv:176:7
					decoded_instr_ack_o[i] = issue_ack_i[i] & ~issue_full[i];
				end
		end
	end
	// Trace: core/scoreboard.sv:182:3
	// removed localparam type ariane_pkg_fu_op
	function automatic ariane_pkg_is_rd_fpr;
		// Trace: core/include/ariane_pkg.sv:597:38
		input reg [7:0] op;
		// Trace: core/include/ariane_pkg.sv:598:5
		(* full_case, parallel_case *)
		case (op)
			8'd96, 8'd97, 8'd98, 8'd99, 8'd104, 8'd105, 8'd106, 8'd107, 8'd108, 8'd109, 8'd110, 8'd111, 8'd112, 8'd113, 8'd115, 8'd116, 8'd117, 8'd119, 8'd122, 8'd123, 8'd124, 8'd125, 8'd126, 8'd133, 8'd134, 8'd135, 8'd136, 8'd183: ariane_pkg_is_rd_fpr = 1'b1;
			default: ariane_pkg_is_rd_fpr = 1'b0;
		endcase
	endfunction
	function automatic [7:0] sv2v_cast_8;
		input reg [7:0] inp;
		sv2v_cast_8 = inp;
	endfunction
	function automatic [((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) - 1:0] sv2v_cast_7EDCF;
		input reg [((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) - 1:0] inp;
		sv2v_cast_7EDCF = inp;
	endfunction
	always @(*) begin : issue_fifo
		if (_sv2v_0)
			;
		// Trace: core/scoreboard.sv:184:5
		mem_n = mem_q;
		// Trace: core/scoreboard.sv:185:5
		num_issue = 1'sb0;
		// Trace: core/scoreboard.sv:188:5
		begin : sv2v_autoblock_3
			// Trace: core/scoreboard.sv:188:10
			reg [31:0] i;
			// Trace: core/scoreboard.sv:188:10
			for (i = 0; i < CVA6Cfg[16841-:32]; i = i + 1)
				begin
					// Trace: core/scoreboard.sv:189:7
					if ((decoded_instr_valid_i[i] && decoded_instr_ack_o[i]) && !flush_unissued_instr_i) begin
						// Trace: core/scoreboard.sv:192:9
						num_issue = num_issue + 'd1;
						// Trace: core/scoreboard.sv:193:9
						mem_n[issue_pointer[(CVA6Cfg[16841-:32] >= 0 ? i : CVA6Cfg[16841-:32] - i) * CVA6Cfg[16503-:32]+:CVA6Cfg[16503-:32]] * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))+:3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))] = {2'b10, CVA6Cfg[16471] && ariane_pkg_is_rd_fpr(decoded_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)]), sv2v_cast_7EDCF(decoded_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 0 : ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) + (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))+:((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))])};
					end
				end
		end
		begin : sv2v_autoblock_4
			// Trace: core/scoreboard.sv:205:10
			reg [31:0] i;
			// Trace: core/scoreboard.sv:205:10
			for (i = 0; i < CVA6Cfg[16535-:32]; i = i + 1)
				begin
					// Trace: core/scoreboard.sv:207:7
					if ((mem_q[(i * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) - 1) - ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) - 1)-:((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] == 4'd0) && mem_q[(i * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + (2 + (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 0))])
						// Trace: core/scoreboard.sv:207:67
						mem_n[(i * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) - 1) - ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : -(4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))] = 1'b1;
				end
		end
		begin : sv2v_autoblock_5
			// Trace: core/scoreboard.sv:213:10
			reg [31:0] i;
			// Trace: core/scoreboard.sv:213:10
			for (i = 0; i < CVA6Cfg[16401-:32]; i = i + 1)
				begin
					// Trace: core/scoreboard.sv:216:7
					if (wt_valid_i[i] && mem_q[(trans_id_i[i * CVA6Cfg[16503-:32]+:CVA6Cfg[16503-:32]] * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + (2 + (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 0))]) begin
						// Trace: core/scoreboard.sv:217:9
						if (mem_q[(trans_id_i[i * CVA6Cfg[16503-:32]+:CVA6Cfg[16503-:32]] * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) - 1) - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 3) : -1)] && mem_q[(trans_id_i[i * CVA6Cfg[16503-:32]+:CVA6Cfg[16503-:32]] * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) - 1) - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 1) : -3)]) begin
							begin
								// Trace: core/scoreboard.sv:218:11
								if (mem_q[(trans_id_i[i * CVA6Cfg[16503-:32]+:CVA6Cfg[16503-:32]] * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) - 1) - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 2) : -2)]) begin
									// Trace: core/scoreboard.sv:219:13
									mem_n[(trans_id_i[i * CVA6Cfg[16503-:32]+:CVA6Cfg[16503-:32]] * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) - 1) - ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : -(4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))] = 1'b1;
									// Trace: core/scoreboard.sv:220:13
									mem_n[((sv2v_cast_8(trans_id_i[i * CVA6Cfg[16503-:32]+:CVA6Cfg[16503-:32]]) - 1) * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) - 1) - ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : -(4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))] = 1'b1;
								end
								else
									// Trace: core/scoreboard.sv:222:13
									mem_n[(trans_id_i[i * CVA6Cfg[16503-:32]+:CVA6Cfg[16503-:32]] * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) - 1) - ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : -(4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))] = 1'b0;
							end
						end
						else
							// Trace: core/scoreboard.sv:225:11
							mem_n[(trans_id_i[i * CVA6Cfg[16503-:32]+:CVA6Cfg[16503-:32]] * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) - 1) - ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : -(4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))] = 1'b1;
						// Trace: core/scoreboard.sv:227:9
						mem_n[(trans_id_i[i * CVA6Cfg[16503-:32]+:CVA6Cfg[16503-:32]] * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) - 1) - ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) >= (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) + 1 : ((4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + 1) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 1)-:((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) >= (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) + 1 : ((4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + 1)] = wbdata_i[i * CVA6Cfg[17102-:32]+:CVA6Cfg[17102-:32]];
						if (CVA6Cfg[1321])
							// Trace: core/scoreboard.sv:230:11
							mem_n[(trans_id_i[i * CVA6Cfg[16503-:32]+:CVA6Cfg[16503-:32]] * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) - 1) - ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4) - (((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) - 1) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] - 1)))) : ((0 + ((((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) - 1) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] - 1)) - ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) - 1)-:scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]] = resolved_branch_i[bp_resolve_t_bp_resolve_t_CVA6Cfg[17070-:32] + 4-:((bp_resolve_t_bp_resolve_t_CVA6Cfg[17070-:32] + 4) >= 5 ? bp_resolve_t_bp_resolve_t_CVA6Cfg[17070-:32] + 0 : 6 - (bp_resolve_t_bp_resolve_t_CVA6Cfg[17070-:32] + 4))];
						if (mem_n[(trans_id_i[i * CVA6Cfg[16503-:32]+:CVA6Cfg[16503-:32]] * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) - 1) - ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) - 1)-:((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] == 4'd9) begin
							begin
								// Trace: core/scoreboard.sv:233:11
								if (x_we_i)
									// Trace: core/scoreboard.sv:233:23
									mem_n[(trans_id_i[i * CVA6Cfg[16503-:32]+:CVA6Cfg[16503-:32]] * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) - 1) - ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) - 1)-:((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = x_rd_i;
								else
									// Trace: core/scoreboard.sv:234:16
									mem_n[(trans_id_i[i * CVA6Cfg[16503-:32]+:CVA6Cfg[16503-:32]] * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) - 1) - ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) - 1)-:((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] = 5'b00000;
							end
						end
						if (ex_i[(i * ((((exception_t_exception_t_CVA6Cfg[17102-:32] + exception_t_exception_t_CVA6Cfg[17102-:32]) + exception_t_exception_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((exception_t_exception_t_CVA6Cfg[17102-:32] + exception_t_exception_t_CVA6Cfg[17102-:32]) + exception_t_exception_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((exception_t_exception_t_CVA6Cfg[17102-:32] + exception_t_exception_t_CVA6Cfg[17102-:32]) + exception_t_exception_t_CVA6Cfg[17006-:32]) + 33))) + ((((exception_t_exception_t_CVA6Cfg[17102-:32] + exception_t_exception_t_CVA6Cfg[17102-:32]) + exception_t_exception_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? 0 : ((exception_t_exception_t_CVA6Cfg[17102-:32] + exception_t_exception_t_CVA6Cfg[17102-:32]) + exception_t_exception_t_CVA6Cfg[17006-:32]) + 33)])
							// Trace: core/scoreboard.sv:237:28
							mem_n[(trans_id_i[i * CVA6Cfg[16503-:32]+:CVA6Cfg[16503-:32]] * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) - 1) - ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) >= ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5) ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) - ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)) + 1 : (((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5) - (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))) + 1) - (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))) - 1)-:((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) >= ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5) ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) - ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)) + 1 : (((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5) - (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))) + 1)] = ex_i[((((exception_t_exception_t_CVA6Cfg[17102-:32] + exception_t_exception_t_CVA6Cfg[17102-:32]) + exception_t_exception_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? 0 : ((exception_t_exception_t_CVA6Cfg[17102-:32] + exception_t_exception_t_CVA6Cfg[17102-:32]) + exception_t_exception_t_CVA6Cfg[17006-:32]) + 33) + (i * ((((exception_t_exception_t_CVA6Cfg[17102-:32] + exception_t_exception_t_CVA6Cfg[17102-:32]) + exception_t_exception_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((exception_t_exception_t_CVA6Cfg[17102-:32] + exception_t_exception_t_CVA6Cfg[17102-:32]) + exception_t_exception_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((exception_t_exception_t_CVA6Cfg[17102-:32] + exception_t_exception_t_CVA6Cfg[17102-:32]) + exception_t_exception_t_CVA6Cfg[17006-:32]) + 33)))+:((((exception_t_exception_t_CVA6Cfg[17102-:32] + exception_t_exception_t_CVA6Cfg[17102-:32]) + exception_t_exception_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((exception_t_exception_t_CVA6Cfg[17102-:32] + exception_t_exception_t_CVA6Cfg[17102-:32]) + exception_t_exception_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((exception_t_exception_t_CVA6Cfg[17102-:32] + exception_t_exception_t_CVA6Cfg[17102-:32]) + exception_t_exception_t_CVA6Cfg[17006-:32]) + 33))];
						else if (CVA6Cfg[16471] && ((mem_q[(trans_id_i[i * CVA6Cfg[16503-:32]+:CVA6Cfg[16503-:32]] * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) - 1) - ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) - 1)-:((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] == 4'd7) || (mem_q[(trans_id_i[i * CVA6Cfg[16503-:32]+:CVA6Cfg[16503-:32]] * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) - 1) - ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) - 1)-:((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] == 4'd8)))
							// Trace: core/scoreboard.sv:240:11
							mem_n[(trans_id_i[i * CVA6Cfg[16503-:32]+:CVA6Cfg[16503-:32]] * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) - 1) - ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) - ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) : ((((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) + ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) + 1)) - 1)) : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) + 1) - ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) - ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) : ((((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) + ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) + 1)) - 1)) - 1)-:((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 34)) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32] + 33)))) + 1)] = ex_i[((((exception_t_exception_t_CVA6Cfg[17102-:32] + exception_t_exception_t_CVA6Cfg[17102-:32]) + exception_t_exception_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? (i * ((((exception_t_exception_t_CVA6Cfg[17102-:32] + exception_t_exception_t_CVA6Cfg[17102-:32]) + exception_t_exception_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((exception_t_exception_t_CVA6Cfg[17102-:32] + exception_t_exception_t_CVA6Cfg[17102-:32]) + exception_t_exception_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((exception_t_exception_t_CVA6Cfg[17102-:32] + exception_t_exception_t_CVA6Cfg[17102-:32]) + exception_t_exception_t_CVA6Cfg[17006-:32]) + 33))) + ((((exception_t_exception_t_CVA6Cfg[17102-:32] + exception_t_exception_t_CVA6Cfg[17102-:32]) + exception_t_exception_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? exception_t_exception_t_CVA6Cfg[17102-:32] + (exception_t_exception_t_CVA6Cfg[17102-:32] + (exception_t_exception_t_CVA6Cfg[17006-:32] + 33)) : (((exception_t_exception_t_CVA6Cfg[17102-:32] + exception_t_exception_t_CVA6Cfg[17102-:32]) + exception_t_exception_t_CVA6Cfg[17006-:32]) + 33) - (exception_t_exception_t_CVA6Cfg[17102-:32] + (exception_t_exception_t_CVA6Cfg[17102-:32] + (exception_t_exception_t_CVA6Cfg[17006-:32] + 33)))) : (((i * ((((exception_t_exception_t_CVA6Cfg[17102-:32] + exception_t_exception_t_CVA6Cfg[17102-:32]) + exception_t_exception_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((exception_t_exception_t_CVA6Cfg[17102-:32] + exception_t_exception_t_CVA6Cfg[17102-:32]) + exception_t_exception_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((exception_t_exception_t_CVA6Cfg[17102-:32] + exception_t_exception_t_CVA6Cfg[17102-:32]) + exception_t_exception_t_CVA6Cfg[17006-:32]) + 33))) + ((((exception_t_exception_t_CVA6Cfg[17102-:32] + exception_t_exception_t_CVA6Cfg[17102-:32]) + exception_t_exception_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? exception_t_exception_t_CVA6Cfg[17102-:32] + (exception_t_exception_t_CVA6Cfg[17102-:32] + (exception_t_exception_t_CVA6Cfg[17006-:32] + 33)) : (((exception_t_exception_t_CVA6Cfg[17102-:32] + exception_t_exception_t_CVA6Cfg[17102-:32]) + exception_t_exception_t_CVA6Cfg[17006-:32]) + 33) - (exception_t_exception_t_CVA6Cfg[17102-:32] + (exception_t_exception_t_CVA6Cfg[17102-:32] + (exception_t_exception_t_CVA6Cfg[17006-:32] + 33))))) + ((exception_t_exception_t_CVA6Cfg[17102-:32] + (exception_t_exception_t_CVA6Cfg[17102-:32] + (exception_t_exception_t_CVA6Cfg[17006-:32] + 33))) >= (exception_t_exception_t_CVA6Cfg[17102-:32] + (exception_t_exception_t_CVA6Cfg[17006-:32] + 34)) ? ((exception_t_exception_t_CVA6Cfg[17102-:32] + (exception_t_exception_t_CVA6Cfg[17102-:32] + (exception_t_exception_t_CVA6Cfg[17006-:32] + 33))) - (exception_t_exception_t_CVA6Cfg[17102-:32] + (exception_t_exception_t_CVA6Cfg[17006-:32] + 34))) + 1 : ((exception_t_exception_t_CVA6Cfg[17102-:32] + (exception_t_exception_t_CVA6Cfg[17006-:32] + 34)) - (exception_t_exception_t_CVA6Cfg[17102-:32] + (exception_t_exception_t_CVA6Cfg[17102-:32] + (exception_t_exception_t_CVA6Cfg[17006-:32] + 33)))) + 1)) - 1)-:((exception_t_exception_t_CVA6Cfg[17102-:32] + (exception_t_exception_t_CVA6Cfg[17102-:32] + (exception_t_exception_t_CVA6Cfg[17006-:32] + 33))) >= (exception_t_exception_t_CVA6Cfg[17102-:32] + (exception_t_exception_t_CVA6Cfg[17006-:32] + 34)) ? ((exception_t_exception_t_CVA6Cfg[17102-:32] + (exception_t_exception_t_CVA6Cfg[17102-:32] + (exception_t_exception_t_CVA6Cfg[17006-:32] + 33))) - (exception_t_exception_t_CVA6Cfg[17102-:32] + (exception_t_exception_t_CVA6Cfg[17006-:32] + 34))) + 1 : ((exception_t_exception_t_CVA6Cfg[17102-:32] + (exception_t_exception_t_CVA6Cfg[17006-:32] + 34)) - (exception_t_exception_t_CVA6Cfg[17102-:32] + (exception_t_exception_t_CVA6Cfg[17102-:32] + (exception_t_exception_t_CVA6Cfg[17006-:32] + 33)))) + 1)];
					end
				end
		end
		if (CVA6Cfg[16809]) begin
			begin
				// Trace: core/scoreboard.sv:249:7
				if (bmiss) begin
					begin
						// Trace: core/scoreboard.sv:250:9
						if (after_flu_wb != issue_pointer[(CVA6Cfg[16841-:32] >= 0 ? 0 : CVA6Cfg[16841-:32]) * CVA6Cfg[16503-:32]+:CVA6Cfg[16503-:32]])
							// Trace: core/scoreboard.sv:251:11
							mem_n[(after_flu_wb * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 1)] = 1'b1;
					end
				end
			end
		end
		begin : sv2v_autoblock_6
			// Trace: core/scoreboard.sv:260:10
			reg signed [31:0] i;
			// Trace: core/scoreboard.sv:260:10
			for (i = 0; i < CVA6Cfg[16873-:32]; i = i + 1)
				begin
					// Trace: core/scoreboard.sv:261:7
					if (commit_ack_i[i]) begin
						// Trace: core/scoreboard.sv:263:9
						mem_n[(commit_pointer_q[i * CVA6Cfg[16503-:32]+:CVA6Cfg[16503-:32]] * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + (2 + (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 0))] = 1'b0;
						// Trace: core/scoreboard.sv:264:9
						mem_n[(commit_pointer_q[i * CVA6Cfg[16503-:32]+:CVA6Cfg[16503-:32]] * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 1)] = 1'b0;
						// Trace: core/scoreboard.sv:265:9
						mem_n[(commit_pointer_q[i * CVA6Cfg[16503-:32]+:CVA6Cfg[16503-:32]] * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) - 1) - ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : -(4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))] = 1'b0;
					end
				end
		end
		if (flush_i)
			// Trace: core/scoreboard.sv:273:7
			begin : sv2v_autoblock_7
				// Trace: core/scoreboard.sv:273:12
				reg [31:0] i;
				// Trace: core/scoreboard.sv:273:12
				for (i = 0; i < CVA6Cfg[16535-:32]; i = i + 1)
					begin
						// Trace: core/scoreboard.sv:275:9
						mem_n[(i * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + (2 + (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 0))] = 1'b0;
						// Trace: core/scoreboard.sv:276:9
						mem_n[(i * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 1)] = 1'b0;
						// Trace: core/scoreboard.sv:277:9
						mem_n[(i * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) - 1) - ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : -(4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))] = 1'b0;
						// Trace: core/scoreboard.sv:278:9
						mem_n[(i * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) - 1) - ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) : (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)) : -((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) : (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))] = 1'b0;
					end
			end
	end
	// Trace: core/scoreboard.sv:283:3
	assign bmiss = resolved_branch_i[1 + (bp_resolve_t_bp_resolve_t_CVA6Cfg[17070-:32] + (bp_resolve_t_bp_resolve_t_CVA6Cfg[17070-:32] + 4))] && resolved_branch_i[4];
	// Trace: core/scoreboard.sv:284:3
	localparam ariane_pkg_FLU_WB = 0;
	assign after_flu_wb = trans_id_i[0+:CVA6Cfg[16503-:32]] + 'd1;
	// Trace: core/scoreboard.sv:287:3
	generate
		if (CVA6Cfg[16873-:32] == 2) begin : gen_commit_ports
			// Trace: core/scoreboard.sv:288:5
			assign num_commit = commit_ack_i[1] + commit_ack_i[0];
		end
		else begin : gen_one_commit_port
			// Trace: core/scoreboard.sv:290:5
			assign num_commit = commit_ack_i[0];
		end
	endgenerate
	// Trace: core/scoreboard.sv:293:3
	assign commit_pointer_n[0+:CVA6Cfg[16503-:32]] = (flush_i ? {CVA6Cfg[16503-:32] * 1 {1'sb0}} : commit_pointer_q[0+:CVA6Cfg[16503-:32]] + num_commit);
	// Trace: core/scoreboard.sv:295:3
	always @(*) begin : assign_issue_pointer_n
		if (_sv2v_0)
			;
		// Trace: core/scoreboard.sv:296:5
		issue_pointer_n = issue_pointer[(CVA6Cfg[16841-:32] >= 0 ? num_issue : CVA6Cfg[16841-:32] - num_issue) * CVA6Cfg[16503-:32]+:CVA6Cfg[16503-:32]];
		// Trace: core/scoreboard.sv:297:5
		if (flush_i)
			// Trace: core/scoreboard.sv:297:18
			issue_pointer_n = 1'sb0;
	end
	// Trace: core/scoreboard.sv:301:3
	genvar _gv_k_5;
	generate
		for (_gv_k_5 = 1; _gv_k_5 < CVA6Cfg[16873-:32]; _gv_k_5 = _gv_k_5 + 1) begin : gen_cnt_incr
			localparam k = _gv_k_5;
			// Trace: core/scoreboard.sv:302:5
			assign commit_pointer_n[k * CVA6Cfg[16503-:32]+:CVA6Cfg[16503-:32]] = (flush_i ? {CVA6Cfg[16503-:32] * 1 {1'sb0}} : commit_pointer_n[0+:CVA6Cfg[16503-:32]] + $unsigned(k));
		end
	endgenerate
	// Trace: core/scoreboard.sv:309:3
	reg [(CVA6Cfg[16535-:32] >= 0 ? (32 * (CVA6Cfg[16535-:32] + 1)) - 1 : (32 * (1 - CVA6Cfg[16535-:32])) + (CVA6Cfg[16535-:32] - 1)):(CVA6Cfg[16535-:32] >= 0 ? 0 : CVA6Cfg[16535-:32] + 0)] gpr_clobber_vld;
	// Trace: core/scoreboard.sv:310:3
	reg [(CVA6Cfg[16535-:32] >= 0 ? (32 * (CVA6Cfg[16535-:32] + 1)) - 1 : (32 * (1 - CVA6Cfg[16535-:32])) + (CVA6Cfg[16535-:32] - 1)):(CVA6Cfg[16535-:32] >= 0 ? 0 : CVA6Cfg[16535-:32] + 0)] fpr_clobber_vld;
	// Trace: core/scoreboard.sv:311:3
	reg [(CVA6Cfg[16535-:32] >= 0 ? ((CVA6Cfg[16535-:32] + 1) * 4) - 1 : ((1 - CVA6Cfg[16535-:32]) * 4) + ((CVA6Cfg[16535-:32] * 4) - 1)):(CVA6Cfg[16535-:32] >= 0 ? 0 : CVA6Cfg[16535-:32] * 4)] clobber_fu;
	// Trace: core/scoreboard.sv:313:3
	always @(*) begin : clobber_assign
		if (_sv2v_0)
			;
		// Trace: core/scoreboard.sv:314:5
		gpr_clobber_vld = 1'sb0;
		// Trace: core/scoreboard.sv:315:5
		fpr_clobber_vld = 1'sb0;
		// Trace: core/scoreboard.sv:318:5
		clobber_fu[(CVA6Cfg[16535-:32] >= 0 ? CVA6Cfg[16535-:32] : CVA6Cfg[16535-:32] - CVA6Cfg[16535-:32]) * 4+:4] = 4'd0;
		// Trace: core/scoreboard.sv:319:5
		begin : sv2v_autoblock_8
			// Trace: core/scoreboard.sv:319:10
			reg [31:0] i;
			// Trace: core/scoreboard.sv:319:10
			for (i = 0; i < 32; i = i + 1)
				begin
					// Trace: core/scoreboard.sv:320:7
					gpr_clobber_vld[(i * (CVA6Cfg[16535-:32] >= 0 ? CVA6Cfg[16535-:32] + 1 : 1 - CVA6Cfg[16535-:32])) + (CVA6Cfg[16535-:32] >= 0 ? CVA6Cfg[16535-:32] : CVA6Cfg[16535-:32] - CVA6Cfg[16535-:32])] = 1'b1;
					// Trace: core/scoreboard.sv:321:7
					fpr_clobber_vld[(i * (CVA6Cfg[16535-:32] >= 0 ? CVA6Cfg[16535-:32] + 1 : 1 - CVA6Cfg[16535-:32])) + (CVA6Cfg[16535-:32] >= 0 ? CVA6Cfg[16535-:32] : CVA6Cfg[16535-:32] - CVA6Cfg[16535-:32])] = 1'b1;
				end
		end
		begin : sv2v_autoblock_9
			// Trace: core/scoreboard.sv:325:10
			reg [31:0] i;
			// Trace: core/scoreboard.sv:325:10
			for (i = 0; i < CVA6Cfg[16535-:32]; i = i + 1)
				begin
					// Trace: core/scoreboard.sv:326:7
					gpr_clobber_vld[(mem_q[(i * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) - 1) - ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) - 1)-:((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] * (CVA6Cfg[16535-:32] >= 0 ? CVA6Cfg[16535-:32] + 1 : 1 - CVA6Cfg[16535-:32])) + (CVA6Cfg[16535-:32] >= 0 ? i : CVA6Cfg[16535-:32] - i)] = still_issued[i] & ~mem_q[(i * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 0)];
					// Trace: core/scoreboard.sv:327:7
					fpr_clobber_vld[(mem_q[(i * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) - 1) - ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) - 1)-:((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] * (CVA6Cfg[16535-:32] >= 0 ? CVA6Cfg[16535-:32] + 1 : 1 - CVA6Cfg[16535-:32])) + (CVA6Cfg[16535-:32] >= 0 ? i : CVA6Cfg[16535-:32] - i)] = still_issued[i] & mem_q[(i * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 0)];
					// Trace: core/scoreboard.sv:328:7
					clobber_fu[(CVA6Cfg[16535-:32] >= 0 ? i : CVA6Cfg[16535-:32] - i) * 4+:4] = mem_q[(i * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) - 1) - ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) - 1)-:((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)];
				end
		end
		// Trace: core/scoreboard.sv:332:5
		gpr_clobber_vld[(CVA6Cfg[16535-:32] >= 0 ? 0 : CVA6Cfg[16535-:32]) + 0+:(CVA6Cfg[16535-:32] >= 0 ? CVA6Cfg[16535-:32] + 1 : 1 - CVA6Cfg[16535-:32])] = 1'sb0;
	end
	// Trace: core/scoreboard.sv:335:3
	genvar _gv_k_6;
	function automatic [31:0] sv2v_cast_32;
		input reg [31:0] inp;
		sv2v_cast_32 = inp;
	endfunction
	generate
		for (_gv_k_6 = 0; _gv_k_6 < 32; _gv_k_6 = _gv_k_6 + 1) begin : gen_sel_clobbers
			localparam k = _gv_k_6;
			// Trace: core/scoreboard.sv:337:5
			localparam [31:0] sv2v_uu_i_sel_gpr_clobbers_NumIn = CVA6Cfg[16535-:32] + 1;
			localparam [31:0] sv2v_uu_i_sel_gpr_clobbers_IdxWidth = (sv2v_uu_i_sel_gpr_clobbers_NumIn > 32'd1 ? $unsigned($clog2(sv2v_uu_i_sel_gpr_clobbers_NumIn)) : 32'd1);
			// removed localparam type sv2v_uu_i_sel_gpr_clobbers_idx_t
			// removed localparam type sv2v_uu_i_sel_gpr_clobbers_rr_i
			localparam [sv2v_cast_32((sv2v_cast_32(CVA6Cfg[16535-:32] + 1) > 32'd1 ? $unsigned($clog2(sv2v_cast_32(CVA6Cfg[16535-:32] + 1))) : 32'd1)) - 1:0] sv2v_uu_i_sel_gpr_clobbers_ext_rr_i_0 = 1'sb0;
			rr_arb_tree_ED597 #(
				.NumIn(CVA6Cfg[16535-:32] + 1),
				.ExtPrio(1'b1),
				.AxiVldRdy(1'b1)
			) i_sel_gpr_clobbers(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.flush_i(1'b0),
				.rr_i(sv2v_uu_i_sel_gpr_clobbers_ext_rr_i_0),
				.req_i(gpr_clobber_vld[(CVA6Cfg[16535-:32] >= 0 ? 0 : CVA6Cfg[16535-:32]) + (k * (CVA6Cfg[16535-:32] >= 0 ? CVA6Cfg[16535-:32] + 1 : 1 - CVA6Cfg[16535-:32]))+:(CVA6Cfg[16535-:32] >= 0 ? CVA6Cfg[16535-:32] + 1 : 1 - CVA6Cfg[16535-:32])]),
				.gnt_o(),
				.data_i(clobber_fu),
				.gnt_i(1'b1),
				.req_o(),
				.data_o(rd_clobber_gpr_o[k * 4+:4]),
				.idx_o()
			);
			if (CVA6Cfg[16471]) begin : genblk1
				// Trace: core/scoreboard.sv:356:7
				localparam [31:0] sv2v_uu_i_sel_fpr_clobbers_NumIn = CVA6Cfg[16535-:32] + 1;
				localparam [31:0] sv2v_uu_i_sel_fpr_clobbers_IdxWidth = (sv2v_uu_i_sel_fpr_clobbers_NumIn > 32'd1 ? $unsigned($clog2(sv2v_uu_i_sel_fpr_clobbers_NumIn)) : 32'd1);
				// removed localparam type sv2v_uu_i_sel_fpr_clobbers_idx_t
				// removed localparam type sv2v_uu_i_sel_fpr_clobbers_rr_i
				localparam [sv2v_cast_32((sv2v_cast_32(CVA6Cfg[16535-:32] + 1) > 32'd1 ? $unsigned($clog2(sv2v_cast_32(CVA6Cfg[16535-:32] + 1))) : 32'd1)) - 1:0] sv2v_uu_i_sel_fpr_clobbers_ext_rr_i_0 = 1'sb0;
				rr_arb_tree_ED597 #(
					.NumIn(CVA6Cfg[16535-:32] + 1),
					.ExtPrio(1'b1),
					.AxiVldRdy(1'b1)
				) i_sel_fpr_clobbers(
					.clk_i(clk_i),
					.rst_ni(rst_ni),
					.flush_i(1'b0),
					.rr_i(sv2v_uu_i_sel_fpr_clobbers_ext_rr_i_0),
					.req_i(fpr_clobber_vld[(CVA6Cfg[16535-:32] >= 0 ? 0 : CVA6Cfg[16535-:32]) + (k * (CVA6Cfg[16535-:32] >= 0 ? CVA6Cfg[16535-:32] + 1 : 1 - CVA6Cfg[16535-:32]))+:(CVA6Cfg[16535-:32] >= 0 ? CVA6Cfg[16535-:32] + 1 : 1 - CVA6Cfg[16535-:32])]),
					.gnt_o(),
					.data_i(clobber_fu),
					.gnt_i(1'b1),
					.req_o(),
					.data_o(rd_clobber_fpr_o[k * 4+:4]),
					.idx_o()
				);
			end
		end
	endgenerate
	// Trace: core/scoreboard.sv:381:3
	wire [(CVA6Cfg[16841-:32] * (CVA6Cfg[16535-:32] + CVA6Cfg[16401-:32])) - 1:0] rs1_fwd_req;
	wire [(CVA6Cfg[16841-:32] * (CVA6Cfg[16535-:32] + CVA6Cfg[16401-:32])) - 1:0] rs2_fwd_req;
	wire [(CVA6Cfg[16841-:32] * (CVA6Cfg[16535-:32] + CVA6Cfg[16401-:32])) - 1:0] rs3_fwd_req;
	// Trace: core/scoreboard.sv:383:3
	wire [((CVA6Cfg[16841-:32] * (CVA6Cfg[16535-:32] + CVA6Cfg[16401-:32])) * CVA6Cfg[17102-:32]) - 1:0] rs_data;
	// Trace: core/scoreboard.sv:384:3
	wire [CVA6Cfg[16841-:32] - 1:0] rs1_valid;
	wire [CVA6Cfg[16841-:32] - 1:0] rs2_valid;
	wire [CVA6Cfg[16841-:32] - 1:0] rs3_valid;
	// Trace: core/scoreboard.sv:387:3
	genvar _gv_i_50;
	function automatic ariane_pkg_is_imm_fpr;
		// Trace: core/include/ariane_pkg.sv:578:39
		input reg [7:0] op;
		// Trace: core/include/ariane_pkg.sv:579:5
		(* full_case, parallel_case *)
		case (op)
			8'd104, 8'd105, 8'd110, 8'd111, 8'd112, 8'd113, 8'd133, 8'd134, 8'd135, 8'd136: ariane_pkg_is_imm_fpr = 1'b1;
			default: ariane_pkg_is_imm_fpr = 1'b0;
		endcase
	endfunction
	function automatic ariane_pkg_is_rs1_fpr;
		// Trace: core/include/ariane_pkg.sv:507:39
		input reg [7:0] op;
		// Trace: core/include/ariane_pkg.sv:508:5
		(* full_case, parallel_case *)
		case (op)
			8'd106, 8'd107, 8'd108, 8'd109, 8'd110, 8'd111, 8'd112, 8'd113, 8'd114, 8'd116, 8'd117, 8'd118, 8'd120, 8'd121, 8'd122, 8'd123, 8'd124, 8'd125, 8'd126, 8'd127, 8'd128, 8'd129, 8'd130, 8'd131, 8'd132, 8'd133, 8'd134, 8'd135, 8'd136, 8'd182: ariane_pkg_is_rs1_fpr = 1'b1;
			default: ariane_pkg_is_rs1_fpr = 1'b0;
		endcase
	endfunction
	function automatic ariane_pkg_is_rs2_fpr;
		// Trace: core/include/ariane_pkg.sv:546:39
		input reg [7:0] op;
		// Trace: core/include/ariane_pkg.sv:547:5
		(* full_case, parallel_case *)
		case (op)
			8'd100, 8'd101, 8'd102, 8'd103, 8'd104, 8'd105, 8'd106, 8'd107, 8'd108, 8'd110, 8'd111, 8'd112, 8'd113, 8'd116, 8'd117, 8'd118, 8'd120, 8'd122, 8'd123, 8'd124, 8'd125, 8'd126: ariane_pkg_is_rs2_fpr = 1'b1;
			default: ariane_pkg_is_rs2_fpr = 1'b0;
		endcase
	endfunction
	localparam cva6_config_pkg_CVA6ConfigXlen = 64;
	localparam riscv_XLEN = cva6_config_pkg_CVA6ConfigXlen;
	generate
		for (_gv_i_50 = 0; _gv_i_50 < CVA6Cfg[16841-:32]; _gv_i_50 = _gv_i_50 + 1) begin : genblk8
			localparam i = _gv_i_50;
			genvar _gv_k_7;
			for (_gv_k_7 = 0; $unsigned(_gv_k_7) < CVA6Cfg[16401-:32]; _gv_k_7 = _gv_k_7 + 1) begin : gen_rs_wb
				localparam k = _gv_k_7;
				// Trace: core/scoreboard.sv:389:7
				assign rs1_fwd_req[(i * (CVA6Cfg[16535-:32] + CVA6Cfg[16401-:32])) + k] = ((((mem_q[(trans_id_i[k * CVA6Cfg[16503-:32]+:CVA6Cfg[16503-:32]] * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) - 1) - ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) - 1)-:((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] == rs1_i[i * 5+:5]) & ~mem_q[(trans_id_i[k * CVA6Cfg[16503-:32]+:CVA6Cfg[16503-:32]] * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 1)]) & wt_valid_i[k]) & ~ex_i[(k * ((((exception_t_exception_t_CVA6Cfg[17102-:32] + exception_t_exception_t_CVA6Cfg[17102-:32]) + exception_t_exception_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((exception_t_exception_t_CVA6Cfg[17102-:32] + exception_t_exception_t_CVA6Cfg[17102-:32]) + exception_t_exception_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((exception_t_exception_t_CVA6Cfg[17102-:32] + exception_t_exception_t_CVA6Cfg[17102-:32]) + exception_t_exception_t_CVA6Cfg[17006-:32]) + 33))) + ((((exception_t_exception_t_CVA6Cfg[17102-:32] + exception_t_exception_t_CVA6Cfg[17102-:32]) + exception_t_exception_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? 0 : ((exception_t_exception_t_CVA6Cfg[17102-:32] + exception_t_exception_t_CVA6Cfg[17102-:32]) + exception_t_exception_t_CVA6Cfg[17006-:32]) + 33)]) & (mem_q[(trans_id_i[k * CVA6Cfg[16503-:32]+:CVA6Cfg[16503-:32]] * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 0)] == (CVA6Cfg[16471] && ariane_pkg_is_rs1_fpr(issue_instr_o[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)])));
				// Trace: core/scoreboard.sv:392:7
				assign rs2_fwd_req[(i * (CVA6Cfg[16535-:32] + CVA6Cfg[16401-:32])) + k] = ((((mem_q[(trans_id_i[k * CVA6Cfg[16503-:32]+:CVA6Cfg[16503-:32]] * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) - 1) - ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) - 1)-:((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] == rs2_i[i * 5+:5]) & ~mem_q[(trans_id_i[k * CVA6Cfg[16503-:32]+:CVA6Cfg[16503-:32]] * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 1)]) & wt_valid_i[k]) & ~ex_i[(k * ((((exception_t_exception_t_CVA6Cfg[17102-:32] + exception_t_exception_t_CVA6Cfg[17102-:32]) + exception_t_exception_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((exception_t_exception_t_CVA6Cfg[17102-:32] + exception_t_exception_t_CVA6Cfg[17102-:32]) + exception_t_exception_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((exception_t_exception_t_CVA6Cfg[17102-:32] + exception_t_exception_t_CVA6Cfg[17102-:32]) + exception_t_exception_t_CVA6Cfg[17006-:32]) + 33))) + ((((exception_t_exception_t_CVA6Cfg[17102-:32] + exception_t_exception_t_CVA6Cfg[17102-:32]) + exception_t_exception_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? 0 : ((exception_t_exception_t_CVA6Cfg[17102-:32] + exception_t_exception_t_CVA6Cfg[17102-:32]) + exception_t_exception_t_CVA6Cfg[17006-:32]) + 33)]) & (mem_q[(trans_id_i[k * CVA6Cfg[16503-:32]+:CVA6Cfg[16503-:32]] * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 0)] == (CVA6Cfg[16471] && ariane_pkg_is_rs2_fpr(issue_instr_o[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)])));
				// Trace: core/scoreboard.sv:395:7
				assign rs3_fwd_req[(i * (CVA6Cfg[16535-:32] + CVA6Cfg[16401-:32])) + k] = ((((mem_q[(trans_id_i[k * CVA6Cfg[16503-:32]+:CVA6Cfg[16503-:32]] * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) - 1) - ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) - 1)-:((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] == rs3_i[i * 5+:5]) & ~mem_q[(trans_id_i[k * CVA6Cfg[16503-:32]+:CVA6Cfg[16503-:32]] * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 1)]) & wt_valid_i[k]) & ~ex_i[(k * ((((exception_t_exception_t_CVA6Cfg[17102-:32] + exception_t_exception_t_CVA6Cfg[17102-:32]) + exception_t_exception_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((exception_t_exception_t_CVA6Cfg[17102-:32] + exception_t_exception_t_CVA6Cfg[17102-:32]) + exception_t_exception_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((exception_t_exception_t_CVA6Cfg[17102-:32] + exception_t_exception_t_CVA6Cfg[17102-:32]) + exception_t_exception_t_CVA6Cfg[17006-:32]) + 33))) + ((((exception_t_exception_t_CVA6Cfg[17102-:32] + exception_t_exception_t_CVA6Cfg[17102-:32]) + exception_t_exception_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? 0 : ((exception_t_exception_t_CVA6Cfg[17102-:32] + exception_t_exception_t_CVA6Cfg[17102-:32]) + exception_t_exception_t_CVA6Cfg[17006-:32]) + 33)]) & (mem_q[(trans_id_i[k * CVA6Cfg[16503-:32]+:CVA6Cfg[16503-:32]] * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 0)] == (CVA6Cfg[16471] && ariane_pkg_is_imm_fpr(issue_instr_o[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)])));
				// Trace: core/scoreboard.sv:398:7
				assign rs_data[((i * (CVA6Cfg[16535-:32] + CVA6Cfg[16401-:32])) + k) * CVA6Cfg[17102-:32]+:CVA6Cfg[17102-:32]] = wbdata_i[k * CVA6Cfg[17102-:32]+:CVA6Cfg[17102-:32]];
			end
			genvar _gv_k_8;
			for (_gv_k_8 = 0; $unsigned(_gv_k_8) < CVA6Cfg[16535-:32]; _gv_k_8 = _gv_k_8 + 1) begin : gen_rs_entries
				localparam k = _gv_k_8;
				// Trace: core/scoreboard.sv:401:7
				assign rs1_fwd_req[(i * (CVA6Cfg[16535-:32] + CVA6Cfg[16401-:32])) + (k + CVA6Cfg[16401-:32])] = (((mem_q[(k * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) - 1) - ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) - 1)-:((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] == rs1_i[i * 5+:5]) & still_issued[k]) & mem_q[(k * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) - 1) - ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : -(4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))]) & (mem_q[(k * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 0)] == (CVA6Cfg[16471] && ariane_pkg_is_rs1_fpr(issue_instr_o[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)])));
				// Trace: core/scoreboard.sv:404:7
				assign rs2_fwd_req[(i * (CVA6Cfg[16535-:32] + CVA6Cfg[16401-:32])) + (k + CVA6Cfg[16401-:32])] = (((mem_q[(k * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) - 1) - ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) - 1)-:((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] == rs2_i[i * 5+:5]) & still_issued[k]) & mem_q[(k * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) - 1) - ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : -(4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))]) & (mem_q[(k * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 0)] == (CVA6Cfg[16471] && ariane_pkg_is_rs2_fpr(issue_instr_o[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)])));
				// Trace: core/scoreboard.sv:407:7
				assign rs3_fwd_req[(i * (CVA6Cfg[16535-:32] + CVA6Cfg[16401-:32])) + (k + CVA6Cfg[16401-:32])] = (((mem_q[(k * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) - 1) - ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) - 1)-:((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] == rs3_i[i * 5+:5]) & still_issued[k]) & mem_q[(k * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) - 1) - ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : -(4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))]) & (mem_q[(k * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + 0)] == (CVA6Cfg[16471] && ariane_pkg_is_imm_fpr(issue_instr_o[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)])));
				// Trace: core/scoreboard.sv:410:7
				assign rs_data[((i * (CVA6Cfg[16535-:32] + CVA6Cfg[16401-:32])) + (k + CVA6Cfg[16401-:32])) * CVA6Cfg[17102-:32]+:CVA6Cfg[17102-:32]] = mem_q[(k * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) - 1) - ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) >= (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) + 1 : ((4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + 1) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 1)-:((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) >= (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) + 1 : ((4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + 1)];
			end
			// Trace: core/scoreboard.sv:414:5
			assign rs1_valid_o[i] = rs1_valid[i] & (|rs1_i[i * 5+:5] | (CVA6Cfg[16471] && ariane_pkg_is_rs1_fpr(issue_instr_o[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)])));
			// Trace: core/scoreboard.sv:417:5
			assign rs2_valid_o[i] = rs2_valid[i] & (|rs2_i[i * 5+:5] | (CVA6Cfg[16471] && ariane_pkg_is_rs2_fpr(issue_instr_o[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)])));
			// Trace: core/scoreboard.sv:420:5
			assign rs3_valid_o[i] = (CVA6Cfg[16433-:32] == 3 ? rs3_valid[i] & (|rs3_i[i * 5+:5] | (CVA6Cfg[16471] && ariane_pkg_is_imm_fpr(issue_instr_o[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)]))) : rs3_valid[i]);
			// Trace: core/scoreboard.sv:426:5
			localparam [31:0] sv2v_uu_i_sel_rs1_NumIn = CVA6Cfg[16535-:32] + CVA6Cfg[16401-:32];
			localparam [31:0] sv2v_uu_i_sel_rs1_IdxWidth = (sv2v_uu_i_sel_rs1_NumIn > 32'd1 ? $unsigned($clog2(sv2v_uu_i_sel_rs1_NumIn)) : 32'd1);
			// removed localparam type sv2v_uu_i_sel_rs1_idx_t
			// removed localparam type sv2v_uu_i_sel_rs1_rr_i
			localparam [sv2v_cast_32((sv2v_cast_32(CVA6Cfg[16535-:32] + CVA6Cfg[16401-:32]) > 32'd1 ? $unsigned($clog2(sv2v_cast_32(CVA6Cfg[16535-:32] + CVA6Cfg[16401-:32]))) : 32'd1)) - 1:0] sv2v_uu_i_sel_rs1_ext_rr_i_0 = 1'sb0;
			rr_arb_tree #(
				.NumIn(CVA6Cfg[16535-:32] + CVA6Cfg[16401-:32]),
				.DataWidth(CVA6Cfg[17102-:32]),
				.ExtPrio(1'b1),
				.AxiVldRdy(1'b1)
			) i_sel_rs1(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.flush_i(1'b0),
				.rr_i(sv2v_uu_i_sel_rs1_ext_rr_i_0),
				.req_i(rs1_fwd_req[i * (CVA6Cfg[16535-:32] + CVA6Cfg[16401-:32])+:CVA6Cfg[16535-:32] + CVA6Cfg[16401-:32]]),
				.gnt_o(),
				.data_i(rs_data[CVA6Cfg[17102-:32] * (i * (CVA6Cfg[16535-:32] + CVA6Cfg[16401-:32]))+:CVA6Cfg[17102-:32] * (CVA6Cfg[16535-:32] + CVA6Cfg[16401-:32])]),
				.gnt_i(1'b1),
				.req_o(rs1_valid[i]),
				.data_o(rs1_o[i * CVA6Cfg[17102-:32]+:CVA6Cfg[17102-:32]]),
				.idx_o()
			);
			// Trace: core/scoreboard.sv:445:5
			localparam [31:0] sv2v_uu_i_sel_rs2_NumIn = CVA6Cfg[16535-:32] + CVA6Cfg[16401-:32];
			localparam [31:0] sv2v_uu_i_sel_rs2_IdxWidth = (sv2v_uu_i_sel_rs2_NumIn > 32'd1 ? $unsigned($clog2(sv2v_uu_i_sel_rs2_NumIn)) : 32'd1);
			// removed localparam type sv2v_uu_i_sel_rs2_idx_t
			// removed localparam type sv2v_uu_i_sel_rs2_rr_i
			localparam [sv2v_cast_32((sv2v_cast_32(CVA6Cfg[16535-:32] + CVA6Cfg[16401-:32]) > 32'd1 ? $unsigned($clog2(sv2v_cast_32(CVA6Cfg[16535-:32] + CVA6Cfg[16401-:32]))) : 32'd1)) - 1:0] sv2v_uu_i_sel_rs2_ext_rr_i_0 = 1'sb0;
			rr_arb_tree #(
				.NumIn(CVA6Cfg[16535-:32] + CVA6Cfg[16401-:32]),
				.DataWidth(CVA6Cfg[17102-:32]),
				.ExtPrio(1'b1),
				.AxiVldRdy(1'b1)
			) i_sel_rs2(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.flush_i(1'b0),
				.rr_i(sv2v_uu_i_sel_rs2_ext_rr_i_0),
				.req_i(rs2_fwd_req[i * (CVA6Cfg[16535-:32] + CVA6Cfg[16401-:32])+:CVA6Cfg[16535-:32] + CVA6Cfg[16401-:32]]),
				.gnt_o(),
				.data_i(rs_data[CVA6Cfg[17102-:32] * (i * (CVA6Cfg[16535-:32] + CVA6Cfg[16401-:32]))+:CVA6Cfg[17102-:32] * (CVA6Cfg[16535-:32] + CVA6Cfg[16401-:32])]),
				.gnt_i(1'b1),
				.req_o(rs2_valid[i]),
				.data_o(rs2_o[i * CVA6Cfg[17102-:32]+:CVA6Cfg[17102-:32]]),
				.idx_o()
			);
			// Trace: core/scoreboard.sv:464:5
			wire [(CVA6Cfg[16841-:32] * CVA6Cfg[17102-:32]) - 1:0] rs3;
			// Trace: core/scoreboard.sv:466:5
			localparam [31:0] sv2v_uu_i_sel_rs3_NumIn = CVA6Cfg[16535-:32] + CVA6Cfg[16401-:32];
			localparam [31:0] sv2v_uu_i_sel_rs3_IdxWidth = (sv2v_uu_i_sel_rs3_NumIn > 32'd1 ? $unsigned($clog2(sv2v_uu_i_sel_rs3_NumIn)) : 32'd1);
			// removed localparam type sv2v_uu_i_sel_rs3_idx_t
			// removed localparam type sv2v_uu_i_sel_rs3_rr_i
			localparam [sv2v_cast_32((sv2v_cast_32(CVA6Cfg[16535-:32] + CVA6Cfg[16401-:32]) > 32'd1 ? $unsigned($clog2(sv2v_cast_32(CVA6Cfg[16535-:32] + CVA6Cfg[16401-:32]))) : 32'd1)) - 1:0] sv2v_uu_i_sel_rs3_ext_rr_i_0 = 1'sb0;
			rr_arb_tree #(
				.NumIn(CVA6Cfg[16535-:32] + CVA6Cfg[16401-:32]),
				.DataWidth(CVA6Cfg[17102-:32]),
				.ExtPrio(1'b1),
				.AxiVldRdy(1'b1)
			) i_sel_rs3(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.flush_i(1'b0),
				.rr_i(sv2v_uu_i_sel_rs3_ext_rr_i_0),
				.req_i(rs3_fwd_req[i * (CVA6Cfg[16535-:32] + CVA6Cfg[16401-:32])+:CVA6Cfg[16535-:32] + CVA6Cfg[16401-:32]]),
				.gnt_o(),
				.data_i(rs_data[CVA6Cfg[17102-:32] * (i * (CVA6Cfg[16535-:32] + CVA6Cfg[16401-:32]))+:CVA6Cfg[17102-:32] * (CVA6Cfg[16535-:32] + CVA6Cfg[16401-:32])]),
				.gnt_i(1'b1),
				.req_o(rs3_valid[i]),
				.data_o(rs3[i * CVA6Cfg[17102-:32]+:CVA6Cfg[17102-:32]]),
				.idx_o()
			);
			if (CVA6Cfg[16433-:32] == 3) begin : gen_gp_three_port
				// Trace: core/scoreboard.sv:486:7
				assign rs3_o[i * (rs3_len_t_CVA6Cfg[16433-:32] == 3 ? rs3_len_t_CVA6Cfg[17102-:32] : rs3_len_t_CVA6Cfg[16469-:32])+:(rs3_len_t_CVA6Cfg[16433-:32] == 3 ? rs3_len_t_CVA6Cfg[17102-:32] : rs3_len_t_CVA6Cfg[16469-:32])] = rs3[(i * CVA6Cfg[17102-:32]) + 63-:64];
			end
			else begin : gen_fp_three_port
				// Trace: core/scoreboard.sv:488:7
				assign rs3_o[i * (rs3_len_t_CVA6Cfg[16433-:32] == 3 ? rs3_len_t_CVA6Cfg[17102-:32] : rs3_len_t_CVA6Cfg[16469-:32])+:(rs3_len_t_CVA6Cfg[16433-:32] == 3 ? rs3_len_t_CVA6Cfg[17102-:32] : rs3_len_t_CVA6Cfg[16469-:32])] = rs3[(i * CVA6Cfg[17102-:32]) + (CVA6Cfg[16469-:32] - 1)-:CVA6Cfg[16469-:32]];
			end
		end
	endgenerate
	// Trace: core/scoreboard.sv:494:3
	function automatic [(3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) - 1:0] sv2v_cast_F037B;
		input reg [(3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) - 1:0] inp;
		sv2v_cast_F037B = inp;
	endfunction
	always @(posedge clk_i or negedge rst_ni) begin : regs
		// Trace: core/scoreboard.sv:495:5
		if (!rst_ni) begin
			// Trace: core/scoreboard.sv:496:7
			mem_q <= {CVA6Cfg[16535-:32] {sv2v_cast_F037B(0)}};
			// Trace: core/scoreboard.sv:497:7
			commit_pointer_q <= 1'sb0;
			// Trace: core/scoreboard.sv:498:7
			issue_pointer_q <= 1'sb0;
		end
		else begin
			// Trace: core/scoreboard.sv:500:7
			issue_pointer_q <= issue_pointer_n;
			// Trace: core/scoreboard.sv:501:7
			mem_q <= mem_n;
			// Trace: core/scoreboard.sv:502:7
			mem_q[(x_id_i * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) - 1) - ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) - 1)-:((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] <= (x_transaction_accepted_i && ~x_issue_writeback_i ? 5'b00000 : mem_n[(x_id_i * (3 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) - 1) - ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) - 1)-:((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)]);
			// Trace: core/scoreboard.sv:503:7
			commit_pointer_q <= commit_pointer_n;
		end
	end
	// Trace: core/scoreboard.sv:508:3
	assign rvfi_issue_pointer_o = issue_pointer[CVA6Cfg[16503-:32] * (CVA6Cfg[16841-:32] >= 0 ? (CVA6Cfg[16841-:32] >= 0 ? (CVA6Cfg[16841-:32] - 1) - (CVA6Cfg[16841-:32] - 1) : CVA6Cfg[16841-:32] - 1) : CVA6Cfg[16841-:32] - (CVA6Cfg[16841-:32] >= 0 ? (CVA6Cfg[16841-:32] - 1) - (CVA6Cfg[16841-:32] - 1) : CVA6Cfg[16841-:32] - 1))+:CVA6Cfg[16503-:32] * CVA6Cfg[16841-:32]];
	// Trace: core/scoreboard.sv:509:3
	assign rvfi_commit_pointer_o = commit_pointer_q;
	// Trace: core/scoreboard.sv:512:3
	// Trace: core/scoreboard.sv:518:3
	// removed an assertion item
	// assert property (@(posedge clk_i) disable iff (!rst_ni)
	// 	rd_clobber_gpr_o[0] == ariane_pkg_NONE
	// ) else begin
	// 	// Trace: core/scoreboard.sv:519:8
	// 	$fatal(1, "RD 0 should not bet set");
	// end
	// Trace: core/scoreboard.sv:521:3
	// removed an assertion item
	// assert property (@(posedge clk_i) disable iff (!rst_ni)
	// 	(commit_ack_i[0] |-> commit_instr_o[0].valid)
	// ) else begin
	// 	// Trace: core/scoreboard.sv:523:8
	// 	$fatal(1, "Commit acknowledged but instruction is not valid");
	// end
	// Trace: core/scoreboard.sv:524:3
	generate
		if (CVA6Cfg[16873-:32] == 2) begin : gen_two_commit_ports
			// Trace: core/scoreboard.sv:525:5
			// removed an assertion item
			// assert property (@(posedge clk_i) disable iff (!rst_ni)
			// 	(commit_ack_i[1] |-> commit_instr_o[1].valid)
			// ) else begin
			// 	// Trace: core/scoreboard.sv:527:10
			// 	$fatal(1, "Commit acknowledged but instruction is not valid");
			// end
		end
	endgenerate
	// Trace: core/scoreboard.sv:530:3
	genvar _gv_i_51;
	generate
		for (_gv_i_51 = 0; _gv_i_51 < CVA6Cfg[16841-:32]; _gv_i_51 = _gv_i_51 + 1) begin : genblk10
			localparam i = _gv_i_51;
			// Trace: core/scoreboard.sv:531:5
			// removed an assertion item
			// assert property (@(posedge clk_i) disable iff (!rst_ni)
			// 	(issue_ack_i[i] |-> issue_instr_valid_o[i])
			// ) else begin
			// 	// Trace: core/scoreboard.sv:533:10
			// 	$fatal(1, "Issue acknowledged but instruction is not valid");
			// end
		end
	endgenerate
	// Trace: core/scoreboard.sv:538:3
	genvar _gv_i_52;
	generate
		for (_gv_i_52 = 0; _gv_i_52 < CVA6Cfg[16401-:32]; _gv_i_52 = _gv_i_52 + 1) begin : genblk11
			localparam i = _gv_i_52;
			genvar _gv_j_5;
			for (_gv_j_5 = 0; _gv_j_5 < CVA6Cfg[16401-:32]; _gv_j_5 = _gv_j_5 + 1) begin : genblk1
				localparam j = _gv_j_5;
				// Trace: core/scoreboard.sv:540:7
				// removed an assertion item
				// assert property (@(posedge clk_i) disable iff (!rst_ni)
				// 	((wt_valid_i[i] && wt_valid_i[j]) && (i != j) |-> trans_id_i[i] != trans_id_i[j])
				// ) else begin
				// 	// Trace: core/scoreboard.sv:543:9
				// 	$fatal(1, "Two or more functional units are retiring instructions with the same transaction id!");
				// end
			end
		end
	endgenerate
	initial _sv2v_0 = 0;
endmodule
