module hpdcache_mem_to_axi_read_9FA2A_A93C0 (
	req_ready_o,
	req_valid_i,
	req_i,
	resp_ready_i,
	resp_valid_o,
	resp_o,
	axi_ar_valid_o,
	axi_ar_o,
	axi_ar_ready_i,
	axi_r_valid_i,
	axi_r_i,
	axi_r_ready_o
);
	// removed localparam type ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_AddrWidth_type
	// removed localparam type ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_IdWidth_type
	// removed localparam type ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth_type
	parameter signed [31:0] ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_AddrWidth = 0;
	parameter signed [31:0] ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_IdWidth = 0;
	parameter signed [31:0] ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth = 0;
	// removed localparam type hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg_type
	parameter [1349:0] hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg = 0;
	// removed localparam type hpdcache_mem_resp_r_t_hpdcache_mem_resp_r_t_HPDcacheCfg_type
	parameter [1349:0] hpdcache_mem_resp_r_t_hpdcache_mem_resp_r_t_HPDcacheCfg = 0;
	// removed localparam type r_chan_t_axi_r_chan_t_axi_r_chan_t_CVA6Cfg_type
	// removed localparam type r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules_type
	parameter [17102:0] r_chan_t_axi_r_chan_t_axi_r_chan_t_CVA6Cfg = 0;
	parameter signed [31:0] r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules = 0;
	reg _sv2v_0;
	// removed import hpdcache_pkg::*;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_read.sv:29:20
	// removed localparam type hpdcache_mem_req_t
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_read.sv:30:20
	// removed localparam type hpdcache_mem_resp_r_t
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_read.sv:31:20
	// removed localparam type ar_chan_t
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_read.sv:32:20
	// removed localparam type r_chan_t
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_read.sv:35:5
	output wire req_ready_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_read.sv:36:5
	input wire req_valid_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_read.sv:37:5
	input wire [((hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[639-:32] + 11) + hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[607-:32]) + 6:0] req_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_read.sv:39:5
	input wire resp_ready_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_read.sv:40:5
	output wire resp_valid_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_read.sv:41:5
	output wire [((2 + hpdcache_mem_resp_r_t_hpdcache_mem_resp_r_t_HPDcacheCfg[607-:32]) + hpdcache_mem_resp_r_t_hpdcache_mem_resp_r_t_HPDcacheCfg[575-:32]) + 0:0] resp_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_read.sv:43:5
	output wire axi_ar_valid_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_read.sv:44:5
	output wire [(((ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_IdWidth + ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_AddrWidth) + 29) + ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth) - 1:0] axi_ar_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_read.sv:45:5
	input wire axi_ar_ready_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_read.sv:47:5
	input wire axi_r_valid_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_read.sv:48:5
	input wire [(((r_chan_t_axi_r_chan_t_axi_r_chan_t_CVA6Cfg[9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + r_chan_t_axi_r_chan_t_axi_r_chan_t_CVA6Cfg[9151 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9151 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9151 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9151 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + 3) + r_chan_t_axi_r_chan_t_axi_r_chan_t_CVA6Cfg[9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) - 1:0] axi_r_i;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_read.sv:49:5
	output wire axi_r_ready_o;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_read.sv:52:5
	wire lock;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_read.sv:53:5
	// removed localparam type axi_pkg_cache_t
	wire [3:0] cache;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_read.sv:54:5
	// removed localparam type hpdcache_pkg_hpdcache_mem_error_e
	reg [1:0] resp;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_read.sv:56:5
	// removed localparam type hpdcache_pkg_hpdcache_mem_command_e
	// removed localparam type hpdcache_pkg_hpdcache_mem_atomic_e
	assign lock = (req_i[6-:2] == 2'b10) && (req_i[4-:4] == 4'b1100);
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_read.sv:59:5
	localparam axi_pkg_CACHE_BUFFERABLE = 4'b0001;
	localparam axi_pkg_CACHE_MODIFIABLE = 4'b0010;
	localparam axi_pkg_CACHE_RD_ALLOC = 4'b0100;
	localparam axi_pkg_CACHE_WR_ALLOC = 4'b1000;
	assign cache = (req_i[0] ? ((axi_pkg_CACHE_BUFFERABLE | axi_pkg_CACHE_MODIFIABLE) | axi_pkg_CACHE_RD_ALLOC) | axi_pkg_CACHE_WR_ALLOC : {4 {1'sb0}});
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_read.sv:65:5
	localparam axi_pkg_RESP_DECERR = 2'b11;
	localparam axi_pkg_RESP_SLVERR = 2'b10;
	always @(*) begin : resp_decode_comb
		if (_sv2v_0)
			;
		// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_read.sv:67:9
		case (axi_r_i[r_chan_t_axi_r_chan_t_axi_r_chan_t_CVA6Cfg[9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 2-:((r_chan_t_axi_r_chan_t_axi_r_chan_t_CVA6Cfg[9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 2) >= (1 + (r_chan_t_axi_r_chan_t_axi_r_chan_t_CVA6Cfg[9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0)) ? ((r_chan_t_axi_r_chan_t_axi_r_chan_t_CVA6Cfg[9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 2) - (1 + (r_chan_t_axi_r_chan_t_axi_r_chan_t_CVA6Cfg[9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0))) + 1 : ((1 + (r_chan_t_axi_r_chan_t_axi_r_chan_t_CVA6Cfg[9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0)) - (r_chan_t_axi_r_chan_t_axi_r_chan_t_CVA6Cfg[9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 2)) + 1)])
			axi_pkg_RESP_SLVERR, axi_pkg_RESP_DECERR:
				// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_read.sv:69:35
				resp = 2'b01;
			default:
				// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_read.sv:70:35
				resp = 2'b00;
		endcase
	end
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_read.sv:74:5
	assign req_ready_o = axi_ar_ready_i;
	assign axi_ar_valid_o = req_valid_i;
	assign axi_ar_o[ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_IdWidth + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_AddrWidth + (21 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 7)))-:((ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_IdWidth + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_AddrWidth + (21 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 7)))) >= (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_AddrWidth + (29 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 0))) ? ((ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_IdWidth + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_AddrWidth + (21 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 7)))) - (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_AddrWidth + (29 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 0)))) + 1 : ((ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_AddrWidth + (29 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 0))) - (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_IdWidth + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_AddrWidth + (21 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 7))))) + 1)] = req_i[hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[607-:32] + 6-:((hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[607-:32] + 6) >= 7 ? hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[607-:32] + 0 : 8 - (hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[607-:32] + 6))];
	assign axi_ar_o[ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_AddrWidth + (21 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 7))-:((ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_AddrWidth + (21 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 7))) >= (29 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 0)) ? ((ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_AddrWidth + (21 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 7))) - (29 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 0))) + 1 : ((29 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 0)) - (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_AddrWidth + (21 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 7)))) + 1)] = req_i[hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[639-:32] + (11 + (hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[607-:32] + 6))-:((hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[639-:32] + (11 + (hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[607-:32] + 6))) >= (11 + (hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[607-:32] + 7)) ? ((hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[639-:32] + (11 + (hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[607-:32] + 6))) - (11 + (hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[607-:32] + 7))) + 1 : ((11 + (hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[607-:32] + 7)) - (hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[639-:32] + (11 + (hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[607-:32] + 6)))) + 1)];
	assign axi_ar_o[21 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 7)-:((21 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 7)) >= (21 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 0)) ? ((21 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 7)) - (21 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 0))) + 1 : ((21 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 0)) - (21 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 7))) + 1)] = req_i[11 + (hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[607-:32] + 6)-:((11 + (hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[607-:32] + 6)) >= (3 + (hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[607-:32] + 7)) ? ((11 + (hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[607-:32] + 6)) - (3 + (hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[607-:32] + 7))) + 1 : ((3 + (hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[607-:32] + 7)) - (11 + (hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[607-:32] + 6))) + 1)];
	assign axi_ar_o[17 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 3)-:((17 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 3)) >= (18 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 0)) ? ((17 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 3)) - (18 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 0))) + 1 : ((18 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 0)) - (17 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 3))) + 1)] = req_i[3 + (hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[607-:32] + 6)-:((3 + (hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[607-:32] + 6)) >= (hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[607-:32] + 7) ? ((3 + (hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[607-:32] + 6)) - (hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[607-:32] + 7)) + 1 : ((hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[607-:32] + 7) - (3 + (hpdcache_mem_req_t_hpdcache_mem_req_t_HPDcacheCfg[607-:32] + 6))) + 1)];
	localparam axi_pkg_BURST_INCR = 2'b01;
	assign axi_ar_o[10 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 7)-:((10 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 7)) >= (16 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 0)) ? ((10 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 7)) - (16 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 0))) + 1 : ((16 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 0)) - (10 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 7))) + 1)] = axi_pkg_BURST_INCR;
	assign axi_ar_o[12 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 3)] = lock;
	assign axi_ar_o[7 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 7)-:((7 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 7)) >= (11 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 0)) ? ((7 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 7)) - (11 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 0))) + 1 : ((11 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 0)) - (7 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 7))) + 1)] = cache;
	assign axi_ar_o[7 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 3)-:((7 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 3)) >= (8 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 0)) ? ((7 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 3)) - (8 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 0))) + 1 : ((8 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 0)) - (7 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 3))) + 1)] = 1'sb0;
	assign axi_ar_o[ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 7-:((ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 7) >= (4 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 0)) ? ((ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 7) - (4 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 0))) + 1 : ((4 + (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 0)) - (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 7)) + 1)] = 1'sb0;
	assign axi_ar_o[ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 3-:((ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 3) >= (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 0) ? ((ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 3) - (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 0)) + 1 : ((ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 0) - (ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth + 3)) + 1)] = 1'sb0;
	assign axi_ar_o[ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth - 1-:ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_axi_ar_chan_t_ariane_axi_UserWidth] = 1'sb0;
	// Trace: core/cache_subsystem/hpdcache/rtl/src/utils/hpdcache_mem_to_axi_read.sv:88:5
	assign axi_r_ready_o = resp_ready_i;
	assign resp_valid_o = axi_r_valid_i;
	assign resp_o[2 + (hpdcache_mem_resp_r_t_hpdcache_mem_resp_r_t_HPDcacheCfg[607-:32] + (hpdcache_mem_resp_r_t_hpdcache_mem_resp_r_t_HPDcacheCfg[575-:32] + 0))-:((2 + (hpdcache_mem_resp_r_t_hpdcache_mem_resp_r_t_HPDcacheCfg[607-:32] + (hpdcache_mem_resp_r_t_hpdcache_mem_resp_r_t_HPDcacheCfg[575-:32] + 0))) >= (hpdcache_mem_resp_r_t_hpdcache_mem_resp_r_t_HPDcacheCfg[607-:32] + (hpdcache_mem_resp_r_t_hpdcache_mem_resp_r_t_HPDcacheCfg[575-:32] + 1)) ? ((2 + (hpdcache_mem_resp_r_t_hpdcache_mem_resp_r_t_HPDcacheCfg[607-:32] + (hpdcache_mem_resp_r_t_hpdcache_mem_resp_r_t_HPDcacheCfg[575-:32] + 0))) - (hpdcache_mem_resp_r_t_hpdcache_mem_resp_r_t_HPDcacheCfg[607-:32] + (hpdcache_mem_resp_r_t_hpdcache_mem_resp_r_t_HPDcacheCfg[575-:32] + 1))) + 1 : ((hpdcache_mem_resp_r_t_hpdcache_mem_resp_r_t_HPDcacheCfg[607-:32] + (hpdcache_mem_resp_r_t_hpdcache_mem_resp_r_t_HPDcacheCfg[575-:32] + 1)) - (2 + (hpdcache_mem_resp_r_t_hpdcache_mem_resp_r_t_HPDcacheCfg[607-:32] + (hpdcache_mem_resp_r_t_hpdcache_mem_resp_r_t_HPDcacheCfg[575-:32] + 0)))) + 1)] = resp;
	assign resp_o[hpdcache_mem_resp_r_t_hpdcache_mem_resp_r_t_HPDcacheCfg[607-:32] + (hpdcache_mem_resp_r_t_hpdcache_mem_resp_r_t_HPDcacheCfg[575-:32] + 0)-:((hpdcache_mem_resp_r_t_hpdcache_mem_resp_r_t_HPDcacheCfg[607-:32] + (hpdcache_mem_resp_r_t_hpdcache_mem_resp_r_t_HPDcacheCfg[575-:32] + 0)) >= (hpdcache_mem_resp_r_t_hpdcache_mem_resp_r_t_HPDcacheCfg[575-:32] + 1) ? ((hpdcache_mem_resp_r_t_hpdcache_mem_resp_r_t_HPDcacheCfg[607-:32] + (hpdcache_mem_resp_r_t_hpdcache_mem_resp_r_t_HPDcacheCfg[575-:32] + 0)) - (hpdcache_mem_resp_r_t_hpdcache_mem_resp_r_t_HPDcacheCfg[575-:32] + 1)) + 1 : ((hpdcache_mem_resp_r_t_hpdcache_mem_resp_r_t_HPDcacheCfg[575-:32] + 1) - (hpdcache_mem_resp_r_t_hpdcache_mem_resp_r_t_HPDcacheCfg[607-:32] + (hpdcache_mem_resp_r_t_hpdcache_mem_resp_r_t_HPDcacheCfg[575-:32] + 0))) + 1)] = axi_r_i[r_chan_t_axi_r_chan_t_axi_r_chan_t_CVA6Cfg[9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (r_chan_t_axi_r_chan_t_axi_r_chan_t_CVA6Cfg[9151 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9151 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9151 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9151 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (r_chan_t_axi_r_chan_t_axi_r_chan_t_CVA6Cfg[9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 2))-:((r_chan_t_axi_r_chan_t_axi_r_chan_t_CVA6Cfg[9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (r_chan_t_axi_r_chan_t_axi_r_chan_t_CVA6Cfg[9151 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9151 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9151 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9151 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (r_chan_t_axi_r_chan_t_axi_r_chan_t_CVA6Cfg[9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 2))) >= (r_chan_t_axi_r_chan_t_axi_r_chan_t_CVA6Cfg[9151 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9151 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9151 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9151 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (3 + (r_chan_t_axi_r_chan_t_axi_r_chan_t_CVA6Cfg[9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0))) ? ((r_chan_t_axi_r_chan_t_axi_r_chan_t_CVA6Cfg[9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (r_chan_t_axi_r_chan_t_axi_r_chan_t_CVA6Cfg[9151 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9151 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9151 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9151 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (r_chan_t_axi_r_chan_t_axi_r_chan_t_CVA6Cfg[9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 2))) - (r_chan_t_axi_r_chan_t_axi_r_chan_t_CVA6Cfg[9151 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9151 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9151 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9151 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (3 + (r_chan_t_axi_r_chan_t_axi_r_chan_t_CVA6Cfg[9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0)))) + 1 : ((r_chan_t_axi_r_chan_t_axi_r_chan_t_CVA6Cfg[9151 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9151 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9151 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9151 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (3 + (r_chan_t_axi_r_chan_t_axi_r_chan_t_CVA6Cfg[9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0))) - (r_chan_t_axi_r_chan_t_axi_r_chan_t_CVA6Cfg[9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (r_chan_t_axi_r_chan_t_axi_r_chan_t_CVA6Cfg[9151 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9151 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9151 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9151 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (r_chan_t_axi_r_chan_t_axi_r_chan_t_CVA6Cfg[9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 2)))) + 1)];
	assign resp_o[hpdcache_mem_resp_r_t_hpdcache_mem_resp_r_t_HPDcacheCfg[575-:32] + 0-:((hpdcache_mem_resp_r_t_hpdcache_mem_resp_r_t_HPDcacheCfg[575-:32] + 0) >= 1 ? hpdcache_mem_resp_r_t_hpdcache_mem_resp_r_t_HPDcacheCfg[575-:32] + 0 : 2 - (hpdcache_mem_resp_r_t_hpdcache_mem_resp_r_t_HPDcacheCfg[575-:32] + 0))] = axi_r_i[r_chan_t_axi_r_chan_t_axi_r_chan_t_CVA6Cfg[9151 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9151 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9151 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9151 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (r_chan_t_axi_r_chan_t_axi_r_chan_t_CVA6Cfg[9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 2)-:((r_chan_t_axi_r_chan_t_axi_r_chan_t_CVA6Cfg[9151 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9151 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9151 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9151 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (r_chan_t_axi_r_chan_t_axi_r_chan_t_CVA6Cfg[9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 2)) >= (3 + (r_chan_t_axi_r_chan_t_axi_r_chan_t_CVA6Cfg[9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0)) ? ((r_chan_t_axi_r_chan_t_axi_r_chan_t_CVA6Cfg[9151 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9151 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9151 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9151 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (r_chan_t_axi_r_chan_t_axi_r_chan_t_CVA6Cfg[9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 2)) - (3 + (r_chan_t_axi_r_chan_t_axi_r_chan_t_CVA6Cfg[9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0))) + 1 : ((3 + (r_chan_t_axi_r_chan_t_axi_r_chan_t_CVA6Cfg[9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0)) - (r_chan_t_axi_r_chan_t_axi_r_chan_t_CVA6Cfg[9151 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9151 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9151 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9119 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9151 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (r_chan_t_axi_r_chan_t_axi_r_chan_t_CVA6Cfg[9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 2))) + 1)];
	assign resp_o[0] = axi_r_i[r_chan_t_axi_r_chan_t_axi_r_chan_t_CVA6Cfg[9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9055 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9087 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + (32 + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + ((r_chan_t_axi_r_chan_t_axi_r_chan_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + 0];
	initial _sv2v_0 = 0;
endmodule
