// removed module with interface ports: apb_to_reg
