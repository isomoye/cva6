module wt_dcache_mem_710D7_EEAC2 (
	clk_i,
	rst_ni,
	rd_tag_i,
	rd_idx_i,
	rd_off_i,
	rd_req_i,
	rd_tag_only_i,
	rd_prio_i,
	rd_ack_o,
	rd_vld_bits_o,
	rd_hit_oh_o,
	rd_data_o,
	rd_user_o,
	wr_cl_vld_i,
	wr_cl_nc_i,
	wr_cl_we_i,
	wr_cl_tag_i,
	wr_cl_idx_i,
	wr_cl_off_i,
	wr_cl_data_i,
	wr_cl_user_i,
	wr_cl_data_be_i,
	wr_vld_bits_i,
	wr_req_i,
	wr_ack_o,
	wr_idx_i,
	wr_off_i,
	wr_data_i,
	wr_user_i,
	wr_data_be_i,
	wbuffer_data_i
);
	// removed localparam type wbuffer_t_CVA6Cfg_type
	// removed localparam type wbuffer_t_config_pkg_NrMaxRules_type
	parameter [17102:0] wbuffer_t_CVA6Cfg = 0;
	parameter signed [31:0] wbuffer_t_config_pkg_NrMaxRules = 0;
	reg _sv2v_0;
	// removed import ariane_pkg::*;
	// removed import wt_cache_pkg::*;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:33:15
	localparam config_pkg_NrMaxRules = 16;
	// removed localparam type config_pkg_cache_type_t
	// removed localparam type config_pkg_noc_type_e
	// removed localparam type config_pkg_vm_mode_t
	// removed localparam type config_pkg_cva6_cfg_t
	localparam [17102:0] config_pkg_cva6_cfg_empty = 17103'd0;
	parameter [17102:0] CVA6Cfg = config_pkg_cva6_cfg_empty;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:34:38
	parameter DCACHE_CL_IDX_WIDTH = 0;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:35:38
	// removed localparam type wbuffer_t
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:36:15
	parameter [31:0] NumPorts = 3;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:38:5
	input wire clk_i;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:39:5
	input wire rst_ni;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:42:5
	input wire [(NumPorts * CVA6Cfg[996-:32]) - 1:0] rd_tag_i;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:43:5
	input wire [(NumPorts * DCACHE_CL_IDX_WIDTH) - 1:0] rd_idx_i;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:44:5
	input wire [(NumPorts * CVA6Cfg[868-:32]) - 1:0] rd_off_i;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:45:5
	input wire [NumPorts - 1:0] rd_req_i;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:46:5
	input wire [NumPorts - 1:0] rd_tag_only_i;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:47:5
	input wire [NumPorts - 1:0] rd_prio_i;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:48:5
	output wire [NumPorts - 1:0] rd_ack_o;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:49:5
	output wire [CVA6Cfg[1092-:32] - 1:0] rd_vld_bits_o;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:50:5
	output wire [CVA6Cfg[1092-:32] - 1:0] rd_hit_oh_o;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:51:5
	output wire [CVA6Cfg[17102-:32] - 1:0] rd_data_o;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:52:5
	output wire [CVA6Cfg[900-:32] - 1:0] rd_user_o;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:55:5
	input wire wr_cl_vld_i;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:56:5
	input wire wr_cl_nc_i;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:57:5
	input wire [CVA6Cfg[1092-:32] - 1:0] wr_cl_we_i;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:58:5
	input wire [CVA6Cfg[996-:32] - 1:0] wr_cl_tag_i;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:59:5
	input wire [DCACHE_CL_IDX_WIDTH - 1:0] wr_cl_idx_i;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:60:5
	input wire [CVA6Cfg[868-:32] - 1:0] wr_cl_off_i;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:61:5
	input wire [CVA6Cfg[964-:32] - 1:0] wr_cl_data_i;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:62:5
	input wire [CVA6Cfg[932-:32] - 1:0] wr_cl_user_i;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:63:5
	input wire [(CVA6Cfg[964-:32] / 8) - 1:0] wr_cl_data_be_i;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:64:5
	input wire [CVA6Cfg[1092-:32] - 1:0] wr_vld_bits_i;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:67:5
	input wire [CVA6Cfg[1092-:32] - 1:0] wr_req_i;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:68:5
	output reg wr_ack_o;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:69:5
	input wire [DCACHE_CL_IDX_WIDTH - 1:0] wr_idx_i;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:70:5
	input wire [CVA6Cfg[868-:32] - 1:0] wr_off_i;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:71:5
	input wire [CVA6Cfg[17102-:32] - 1:0] wr_data_i;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:72:5
	input wire [CVA6Cfg[900-:32] - 1:0] wr_user_i;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:73:5
	input wire [(CVA6Cfg[17102-:32] / 8) - 1:0] wr_data_be_i;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:76:5
	input wire [(CVA6Cfg[740-:32] * ((((((((wbuffer_t_CVA6Cfg[996-:32] + (wbuffer_t_CVA6Cfg[1028-:32] - wbuffer_t_CVA6Cfg[9411 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9411 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9379 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9411 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9379 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9379 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9411 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)])) + wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + wbuffer_t_CVA6Cfg[900-:32]) + (wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8)) + (wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8)) + (wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8)) + 1) + wbuffer_t_CVA6Cfg[1092-:32])) - 1:0] wbuffer_data_i;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:79:3
	localparam DCACHE_NUM_BANKS = CVA6Cfg[964-:32] / CVA6Cfg[17102-:32];
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:80:3
	localparam DCACHE_NUM_BANKS_WIDTH = $clog2(DCACHE_NUM_BANKS);
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:83:3
	function automatic [DCACHE_NUM_BANKS - 1:0] dcache_cl_bin2oh;
		// Trace: core/cache_subsystem/wt_dcache_mem.sv:84:7
		input reg [DCACHE_NUM_BANKS_WIDTH - 1:0] in;
		// Trace: core/cache_subsystem/wt_dcache_mem.sv:85:5
		reg [DCACHE_NUM_BANKS - 1:0] out;
		begin
			// Trace: core/cache_subsystem/wt_dcache_mem.sv:86:5
			out = 1'sb0;
			// Trace: core/cache_subsystem/wt_dcache_mem.sv:87:5
			out[in] = 1'b1;
			// Trace: core/cache_subsystem/wt_dcache_mem.sv:88:5
			dcache_cl_bin2oh = out;
		end
	endfunction
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:93:3
	localparam AXI_OFFSET_WIDTH = (CVA6Cfg[16712-:32] == CVA6Cfg[17102-:32] ? $clog2(CVA6Cfg[16712-:32] / 8) + 1 : $clog2(CVA6Cfg[16712-:32] / 8));
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:99:3
	reg [DCACHE_NUM_BANKS - 1:0] bank_req;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:100:3
	reg [DCACHE_NUM_BANKS - 1:0] bank_we;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:101:3
	wire [((DCACHE_NUM_BANKS * CVA6Cfg[1092-:32]) * (CVA6Cfg[17102-:32] / 8)) - 1:0] bank_be;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:102:3
	reg [(DCACHE_NUM_BANKS * DCACHE_CL_IDX_WIDTH) - 1:0] bank_idx;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:103:3
	wire [DCACHE_CL_IDX_WIDTH - 1:0] bank_idx_d;
	reg [DCACHE_CL_IDX_WIDTH - 1:0] bank_idx_q;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:104:3
	wire [CVA6Cfg[868-:32] - 1:0] bank_off_d;
	reg [CVA6Cfg[868-:32] - 1:0] bank_off_q;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:106:3
	wire [((DCACHE_NUM_BANKS * CVA6Cfg[1092-:32]) * CVA6Cfg[17102-:32]) - 1:0] bank_wdata;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:107:3
	wire [((DCACHE_NUM_BANKS * CVA6Cfg[1092-:32]) * CVA6Cfg[17102-:32]) - 1:0] bank_rdata;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:108:3
	wire [(CVA6Cfg[1092-:32] * CVA6Cfg[17102-:32]) - 1:0] rdata_cl;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:109:3
	wire [((DCACHE_NUM_BANKS * CVA6Cfg[1092-:32]) * CVA6Cfg[900-:32]) - 1:0] bank_wuser;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:110:3
	wire [((DCACHE_NUM_BANKS * CVA6Cfg[1092-:32]) * CVA6Cfg[900-:32]) - 1:0] bank_ruser;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:111:3
	wire [(CVA6Cfg[1092-:32] * CVA6Cfg[900-:32]) - 1:0] ruser_cl;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:113:3
	wire [CVA6Cfg[996-:32] - 1:0] rd_tag;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:114:3
	wire [CVA6Cfg[1092-:32] - 1:0] vld_req;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:115:3
	reg vld_we;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:116:3
	wire [CVA6Cfg[1092-:32] - 1:0] vld_wdata;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:117:3
	wire [(CVA6Cfg[1092-:32] * CVA6Cfg[996-:32]) - 1:0] tag_rdata;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:118:3
	wire [DCACHE_CL_IDX_WIDTH - 1:0] vld_addr;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:120:3
	wire [$clog2(NumPorts) - 1:0] vld_sel_d;
	reg [$clog2(NumPorts) - 1:0] vld_sel_q;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:122:3
	wire [CVA6Cfg[740-:32] - 1:0] wbuffer_hit_oh;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:123:3
	wire [(CVA6Cfg[17102-:32] / 8) - 1:0] wbuffer_be;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:124:3
	wire [CVA6Cfg[17102-:32] - 1:0] wbuffer_rdata;
	reg [CVA6Cfg[17102-:32] - 1:0] rdata;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:125:3
	wire [CVA6Cfg[900-:32] - 1:0] wbuffer_ruser;
	reg [CVA6Cfg[900-:32] - 1:0] ruser;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:126:3
	wire [CVA6Cfg[17038-:32] - 1:0] wbuffer_cmp_addr;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:128:3
	wire cmp_en_d;
	reg cmp_en_q;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:129:3
	wire rd_acked;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:130:3
	reg [NumPorts - 1:0] bank_collision;
	wire [NumPorts - 1:0] rd_req_masked;
	wire [NumPorts - 1:0] rd_req_prio;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:144:3
	genvar _gv_k_9;
	generate
		for (_gv_k_9 = 0; _gv_k_9 < DCACHE_NUM_BANKS; _gv_k_9 = _gv_k_9 + 1) begin : gen_bank
			localparam k = _gv_k_9;
			genvar _gv_j_6;
			for (_gv_j_6 = 0; _gv_j_6 < CVA6Cfg[1092-:32]; _gv_j_6 = _gv_j_6 + 1) begin : gen_bank_way
				localparam j = _gv_j_6;
				// Trace: core/cache_subsystem/wt_dcache_mem.sv:146:7
				assign bank_be[((k * CVA6Cfg[1092-:32]) + j) * (CVA6Cfg[17102-:32] / 8)+:CVA6Cfg[17102-:32] / 8] = (wr_cl_we_i[j] & wr_cl_vld_i ? wr_cl_data_be_i[k * (CVA6Cfg[17102-:32] / 8)+:CVA6Cfg[17102-:32] / 8] : (wr_req_i[j] & wr_ack_o ? wr_data_be_i : {CVA6Cfg[17102-:32] / 8 {1'sb0}}));
				// Trace: core/cache_subsystem/wt_dcache_mem.sv:149:7
				assign bank_wdata[((k * CVA6Cfg[1092-:32]) + j) * CVA6Cfg[17102-:32]+:CVA6Cfg[17102-:32]] = (wr_cl_we_i[j] & wr_cl_vld_i ? wr_cl_data_i[k * CVA6Cfg[17102-:32]+:CVA6Cfg[17102-:32]] : wr_data_i);
				// Trace: core/cache_subsystem/wt_dcache_mem.sv:151:7
				assign bank_wuser[((k * CVA6Cfg[1092-:32]) + j) * CVA6Cfg[900-:32]+:CVA6Cfg[900-:32]] = (wr_cl_we_i[j] & wr_cl_vld_i ? wr_cl_user_i[k * CVA6Cfg[900-:32]+:CVA6Cfg[900-:32]] : wr_user_i);
			end
		end
	endgenerate
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:156:3
	assign vld_wdata = wr_vld_bits_i;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:157:3
	assign vld_addr = (wr_cl_vld_i ? wr_cl_idx_i : rd_idx_i[vld_sel_d * DCACHE_CL_IDX_WIDTH+:DCACHE_CL_IDX_WIDTH]);
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:158:3
	assign rd_tag = rd_tag_i[vld_sel_q * CVA6Cfg[996-:32]+:CVA6Cfg[996-:32]];
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:159:3
	assign bank_off_d = (wr_cl_vld_i ? wr_cl_off_i : rd_off_i[vld_sel_d * CVA6Cfg[868-:32]+:CVA6Cfg[868-:32]]);
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:160:3
	assign bank_idx_d = (wr_cl_vld_i ? wr_cl_idx_i : rd_idx_i[vld_sel_d * DCACHE_CL_IDX_WIDTH+:DCACHE_CL_IDX_WIDTH]);
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:161:3
	assign vld_req = (wr_cl_vld_i ? wr_cl_we_i : (rd_acked ? {CVA6Cfg[1092-:32] {1'sb1}} : {CVA6Cfg[1092-:32] {1'sb0}}));
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:166:3
	assign rd_req_prio = rd_req_i & rd_prio_i;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:167:3
	assign rd_req_masked = (|rd_req_prio ? rd_req_prio : rd_req_i);
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:169:3
	wire rd_req;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:170:3
	// removed localparam type sv2v_uu_i_rr_arb_tree_flush_i
	localparam [0:0] sv2v_uu_i_rr_arb_tree_ext_flush_i_0 = 1'sb0;
	localparam [31:0] sv2v_uu_i_rr_arb_tree_NumIn = NumPorts;
	localparam [31:0] sv2v_uu_i_rr_arb_tree_IdxWidth = (sv2v_uu_i_rr_arb_tree_NumIn > 32'd1 ? $unsigned($clog2(sv2v_uu_i_rr_arb_tree_NumIn)) : 32'd1);
	// removed localparam type sv2v_uu_i_rr_arb_tree_idx_t
	// removed localparam type sv2v_uu_i_rr_arb_tree_rr_i
	localparam [sv2v_uu_i_rr_arb_tree_IdxWidth - 1:0] sv2v_uu_i_rr_arb_tree_ext_rr_i_0 = 1'sb0;
	localparam [31:0] sv2v_uu_i_rr_arb_tree_DataWidth = 1;
	// removed localparam type sv2v_uu_i_rr_arb_tree_DataType
	// removed localparam type sv2v_uu_i_rr_arb_tree_data_i
	localparam [(sv2v_uu_i_rr_arb_tree_NumIn * sv2v_uu_i_rr_arb_tree_DataWidth) - 1:0] sv2v_uu_i_rr_arb_tree_ext_data_i_0 = 1'sb0;
	rr_arb_tree #(
		.NumIn(NumPorts),
		.DataWidth(1)
	) i_rr_arb_tree(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(sv2v_uu_i_rr_arb_tree_ext_flush_i_0),
		.rr_i(sv2v_uu_i_rr_arb_tree_ext_rr_i_0),
		.req_i(rd_req_masked),
		.gnt_o(rd_ack_o),
		.data_i(sv2v_uu_i_rr_arb_tree_ext_data_i_0),
		.gnt_i(~wr_cl_vld_i),
		.req_o(rd_req),
		.data_o(),
		.idx_o(vld_sel_d)
	);
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:187:3
	assign rd_acked = rd_req & ~wr_cl_vld_i;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:189:3
	function automatic [DCACHE_CL_IDX_WIDTH - 1:0] sv2v_cast_E965D;
		input reg [DCACHE_CL_IDX_WIDTH - 1:0] inp;
		sv2v_cast_E965D = inp;
	endfunction
	always @(*) begin : p_bank_req
		if (_sv2v_0)
			;
		// Trace: core/cache_subsystem/wt_dcache_mem.sv:190:5
		vld_we = wr_cl_vld_i;
		// Trace: core/cache_subsystem/wt_dcache_mem.sv:191:5
		bank_req = 1'sb0;
		// Trace: core/cache_subsystem/wt_dcache_mem.sv:192:5
		wr_ack_o = 1'sb0;
		// Trace: core/cache_subsystem/wt_dcache_mem.sv:193:5
		bank_we = 1'sb0;
		// Trace: core/cache_subsystem/wt_dcache_mem.sv:194:5
		bank_idx = {DCACHE_NUM_BANKS {sv2v_cast_E965D(wr_idx_i)}};
		// Trace: core/cache_subsystem/wt_dcache_mem.sv:196:5
		begin : sv2v_autoblock_1
			// Trace: core/cache_subsystem/wt_dcache_mem.sv:196:10
			reg signed [31:0] k;
			// Trace: core/cache_subsystem/wt_dcache_mem.sv:196:10
			for (k = 0; k < NumPorts; k = k + 1)
				begin
					// Trace: core/cache_subsystem/wt_dcache_mem.sv:197:7
					bank_collision[k] = rd_off_i[(k * CVA6Cfg[868-:32]) + ((CVA6Cfg[868-:32] - 1) >= CVA6Cfg[16972-:32] ? CVA6Cfg[868-:32] - 1 : ((CVA6Cfg[868-:32] - 1) + ((CVA6Cfg[868-:32] - 1) >= CVA6Cfg[16972-:32] ? ((CVA6Cfg[868-:32] - 1) - CVA6Cfg[16972-:32]) + 1 : (CVA6Cfg[16972-:32] - (CVA6Cfg[868-:32] - 1)) + 1)) - 1)-:((CVA6Cfg[868-:32] - 1) >= CVA6Cfg[16972-:32] ? ((CVA6Cfg[868-:32] - 1) - CVA6Cfg[16972-:32]) + 1 : (CVA6Cfg[16972-:32] - (CVA6Cfg[868-:32] - 1)) + 1)] == wr_off_i[CVA6Cfg[868-:32] - 1:CVA6Cfg[16972-:32]];
				end
		end
		if (wr_cl_vld_i & |wr_cl_we_i) begin
			// Trace: core/cache_subsystem/wt_dcache_mem.sv:201:7
			bank_req = 1'sb1;
			// Trace: core/cache_subsystem/wt_dcache_mem.sv:202:7
			bank_we = 1'sb1;
			// Trace: core/cache_subsystem/wt_dcache_mem.sv:203:7
			bank_idx = {DCACHE_NUM_BANKS {sv2v_cast_E965D(wr_cl_idx_i)}};
		end
		else begin
			// Trace: core/cache_subsystem/wt_dcache_mem.sv:205:7
			if (rd_acked) begin
				begin
					// Trace: core/cache_subsystem/wt_dcache_mem.sv:206:9
					if (!rd_tag_only_i[vld_sel_d]) begin
						// Trace: core/cache_subsystem/wt_dcache_mem.sv:207:11
						bank_req = dcache_cl_bin2oh(rd_off_i[(vld_sel_d * CVA6Cfg[868-:32]) + ((CVA6Cfg[868-:32] - 1) >= CVA6Cfg[16972-:32] ? CVA6Cfg[868-:32] - 1 : ((CVA6Cfg[868-:32] - 1) + ((CVA6Cfg[868-:32] - 1) >= CVA6Cfg[16972-:32] ? ((CVA6Cfg[868-:32] - 1) - CVA6Cfg[16972-:32]) + 1 : (CVA6Cfg[16972-:32] - (CVA6Cfg[868-:32] - 1)) + 1)) - 1)-:((CVA6Cfg[868-:32] - 1) >= CVA6Cfg[16972-:32] ? ((CVA6Cfg[868-:32] - 1) - CVA6Cfg[16972-:32]) + 1 : (CVA6Cfg[16972-:32] - (CVA6Cfg[868-:32] - 1)) + 1)]);
						// Trace: core/cache_subsystem/wt_dcache_mem.sv:209:11
						bank_idx[rd_off_i[(vld_sel_d * CVA6Cfg[868-:32]) + ((CVA6Cfg[868-:32] - 1) >= CVA6Cfg[16972-:32] ? CVA6Cfg[868-:32] - 1 : ((CVA6Cfg[868-:32] - 1) + ((CVA6Cfg[868-:32] - 1) >= CVA6Cfg[16972-:32] ? ((CVA6Cfg[868-:32] - 1) - CVA6Cfg[16972-:32]) + 1 : (CVA6Cfg[16972-:32] - (CVA6Cfg[868-:32] - 1)) + 1)) - 1)-:((CVA6Cfg[868-:32] - 1) >= CVA6Cfg[16972-:32] ? ((CVA6Cfg[868-:32] - 1) - CVA6Cfg[16972-:32]) + 1 : (CVA6Cfg[16972-:32] - (CVA6Cfg[868-:32] - 1)) + 1)] * DCACHE_CL_IDX_WIDTH+:DCACHE_CL_IDX_WIDTH] = rd_idx_i[vld_sel_d * DCACHE_CL_IDX_WIDTH+:DCACHE_CL_IDX_WIDTH];
					end
				end
			end
			if (|wr_req_i) begin
				begin
					// Trace: core/cache_subsystem/wt_dcache_mem.sv:214:9
					if (rd_tag_only_i[vld_sel_d] || !(rd_ack_o[vld_sel_d] && bank_collision[vld_sel_d])) begin
						// Trace: core/cache_subsystem/wt_dcache_mem.sv:215:11
						wr_ack_o = 1'b1;
						// Trace: core/cache_subsystem/wt_dcache_mem.sv:216:11
						bank_req = bank_req | dcache_cl_bin2oh(wr_off_i[CVA6Cfg[868-:32] - 1:CVA6Cfg[16972-:32]]);
						// Trace: core/cache_subsystem/wt_dcache_mem.sv:219:11
						bank_we = dcache_cl_bin2oh(wr_off_i[CVA6Cfg[868-:32] - 1:CVA6Cfg[16972-:32]]);
					end
				end
			end
		end
	end
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:230:3
	wire [(CVA6Cfg[868-:32] - CVA6Cfg[16972-:32]) - 1:0] wr_cl_off;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:231:3
	wire [(CVA6Cfg[868-:32] - CVA6Cfg[16972-:32]) - 1:0] wr_cl_nc_off;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:232:3
	wire [$clog2(CVA6Cfg[740-:32]) - 1:0] wbuffer_hit_idx;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:233:3
	wire [$clog2(CVA6Cfg[1092-:32]) - 1:0] rd_hit_idx;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:235:3
	assign cmp_en_d = |vld_req & ~vld_we;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:238:3
	assign wbuffer_cmp_addr = (wr_cl_vld_i ? {wr_cl_tag_i, wr_cl_idx_i, wr_cl_off_i} : {rd_tag, bank_idx_q, bank_off_q});
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:241:3
	genvar _gv_i_69;
	generate
		for (_gv_i_69 = 0; _gv_i_69 < CVA6Cfg[1092-:32]; _gv_i_69 = _gv_i_69 + 1) begin : gen_tag_cmpsel
			localparam i = _gv_i_69;
			// Trace: core/cache_subsystem/wt_dcache_mem.sv:243:5
			assign rd_hit_oh_o[i] = ((rd_tag == tag_rdata[i * CVA6Cfg[996-:32]+:CVA6Cfg[996-:32]]) & rd_vld_bits_o[i]) & cmp_en_q;
			// Trace: core/cache_subsystem/wt_dcache_mem.sv:245:5
			assign rdata_cl[i * CVA6Cfg[17102-:32]+:CVA6Cfg[17102-:32]] = bank_rdata[((bank_off_q[CVA6Cfg[868-:32] - 1:CVA6Cfg[16972-:32]] * CVA6Cfg[1092-:32]) + i) * CVA6Cfg[17102-:32]+:CVA6Cfg[17102-:32]];
			// Trace: core/cache_subsystem/wt_dcache_mem.sv:246:5
			assign ruser_cl[i * CVA6Cfg[900-:32]+:CVA6Cfg[900-:32]] = bank_ruser[((bank_off_q[CVA6Cfg[868-:32] - 1:CVA6Cfg[16972-:32]] * CVA6Cfg[1092-:32]) + i) * CVA6Cfg[900-:32]+:CVA6Cfg[900-:32]];
		end
	endgenerate
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:249:3
	genvar _gv_k_10;
	generate
		for (_gv_k_10 = 0; _gv_k_10 < CVA6Cfg[740-:32]; _gv_k_10 = _gv_k_10 + 1) begin : gen_wbuffer_hit
			localparam k = _gv_k_10;
			// Trace: core/cache_subsystem/wt_dcache_mem.sv:250:5
			assign wbuffer_hit_oh[k] = |wbuffer_data_i[(k * ((((((((wbuffer_t_CVA6Cfg[996-:32] + (wbuffer_t_CVA6Cfg[1028-:32] - wbuffer_t_CVA6Cfg[9411 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9411 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9379 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9411 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9379 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9379 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9411 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)])) + wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + wbuffer_t_CVA6Cfg[900-:32]) + (wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8)) + (wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8)) + (wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8)) + 1) + wbuffer_t_CVA6Cfg[1092-:32])) + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + (wbuffer_t_CVA6Cfg[1092-:32] + 0)))-:(((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + (wbuffer_t_CVA6Cfg[1092-:32] + 0))) >= ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + (1 + (wbuffer_t_CVA6Cfg[1092-:32] + 0))) ? (((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + (wbuffer_t_CVA6Cfg[1092-:32] + 0))) - ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + (1 + (wbuffer_t_CVA6Cfg[1092-:32] + 0)))) + 1 : (((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + (1 + (wbuffer_t_CVA6Cfg[1092-:32] + 0))) - ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + (wbuffer_t_CVA6Cfg[1092-:32] + 0)))) + 1)] & ({{CVA6Cfg[16972-:32] {1'b0}}, wbuffer_data_i[(k * ((((((((wbuffer_t_CVA6Cfg[996-:32] + (wbuffer_t_CVA6Cfg[1028-:32] - wbuffer_t_CVA6Cfg[9411 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9411 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9379 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9411 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9379 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9379 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9411 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)])) + wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + wbuffer_t_CVA6Cfg[900-:32]) + (wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8)) + (wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8)) + (wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8)) + 1) + wbuffer_t_CVA6Cfg[1092-:32])) + ((wbuffer_t_CVA6Cfg[996-:32] + (wbuffer_t_CVA6Cfg[1028-:32] - wbuffer_t_CVA6Cfg[9411 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9411 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9379 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9411 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9379 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9379 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9411 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)])) + (wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (wbuffer_t_CVA6Cfg[900-:32] + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + (wbuffer_t_CVA6Cfg[1092-:32] + 0)))))))-:(((wbuffer_t_CVA6Cfg[996-:32] + (wbuffer_t_CVA6Cfg[1028-:32] - wbuffer_t_CVA6Cfg[9411 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9411 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9379 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9411 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9379 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9379 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9411 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)])) + (wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (wbuffer_t_CVA6Cfg[900-:32] + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + (wbuffer_t_CVA6Cfg[1092-:32] + 0))))))) >= (wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (wbuffer_t_CVA6Cfg[900-:32] + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + (1 + (wbuffer_t_CVA6Cfg[1092-:32] + 0))))))) ? (((wbuffer_t_CVA6Cfg[996-:32] + (wbuffer_t_CVA6Cfg[1028-:32] - wbuffer_t_CVA6Cfg[9411 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9411 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9379 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9411 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9379 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9379 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9411 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)])) + (wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (wbuffer_t_CVA6Cfg[900-:32] + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + (wbuffer_t_CVA6Cfg[1092-:32] + 0))))))) - (wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (wbuffer_t_CVA6Cfg[900-:32] + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + (1 + (wbuffer_t_CVA6Cfg[1092-:32] + 0)))))))) + 1 : ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (wbuffer_t_CVA6Cfg[900-:32] + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + (1 + (wbuffer_t_CVA6Cfg[1092-:32] + 0))))))) - ((wbuffer_t_CVA6Cfg[996-:32] + (wbuffer_t_CVA6Cfg[1028-:32] - wbuffer_t_CVA6Cfg[9411 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9411 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9379 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9411 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9379 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9379 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9411 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)])) + (wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (wbuffer_t_CVA6Cfg[900-:32] + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + (wbuffer_t_CVA6Cfg[1092-:32] + 0)))))))) + 1)]} == (wbuffer_cmp_addr >> CVA6Cfg[16972-:32]));
		end
	endgenerate
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:253:3
	lzc #(.WIDTH(CVA6Cfg[740-:32])) i_lzc_wbuffer_hit(
		.in_i(wbuffer_hit_oh),
		.cnt_o(wbuffer_hit_idx),
		.empty_o()
	);
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:261:3
	lzc #(.WIDTH(CVA6Cfg[1092-:32])) i_lzc_rd_hit(
		.in_i(rd_hit_oh_o),
		.cnt_o(rd_hit_idx),
		.empty_o()
	);
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:269:3
	assign wbuffer_rdata = wbuffer_data_i[(wbuffer_hit_idx * ((((((((wbuffer_t_CVA6Cfg[996-:32] + (wbuffer_t_CVA6Cfg[1028-:32] - wbuffer_t_CVA6Cfg[9411 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9411 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9379 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9411 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9379 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9379 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9411 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)])) + wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + wbuffer_t_CVA6Cfg[900-:32]) + (wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8)) + (wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8)) + (wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8)) + 1) + wbuffer_t_CVA6Cfg[1092-:32])) + (wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (wbuffer_t_CVA6Cfg[900-:32] + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + (wbuffer_t_CVA6Cfg[1092-:32] + 0))))))-:((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (wbuffer_t_CVA6Cfg[900-:32] + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + (wbuffer_t_CVA6Cfg[1092-:32] + 0)))))) >= (wbuffer_t_CVA6Cfg[900-:32] + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + (1 + (wbuffer_t_CVA6Cfg[1092-:32] + 0)))))) ? ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (wbuffer_t_CVA6Cfg[900-:32] + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + (wbuffer_t_CVA6Cfg[1092-:32] + 0)))))) - (wbuffer_t_CVA6Cfg[900-:32] + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + (1 + (wbuffer_t_CVA6Cfg[1092-:32] + 0))))))) + 1 : ((wbuffer_t_CVA6Cfg[900-:32] + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + (1 + (wbuffer_t_CVA6Cfg[1092-:32] + 0)))))) - (wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] + (wbuffer_t_CVA6Cfg[900-:32] + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + (wbuffer_t_CVA6Cfg[1092-:32] + 0))))))) + 1)];
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:270:3
	assign wbuffer_ruser = wbuffer_data_i[(wbuffer_hit_idx * ((((((((wbuffer_t_CVA6Cfg[996-:32] + (wbuffer_t_CVA6Cfg[1028-:32] - wbuffer_t_CVA6Cfg[9411 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9411 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9379 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9411 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9379 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9379 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9411 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)])) + wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + wbuffer_t_CVA6Cfg[900-:32]) + (wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8)) + (wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8)) + (wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8)) + 1) + wbuffer_t_CVA6Cfg[1092-:32])) + (wbuffer_t_CVA6Cfg[900-:32] + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + (wbuffer_t_CVA6Cfg[1092-:32] + 0)))))-:((wbuffer_t_CVA6Cfg[900-:32] + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + (wbuffer_t_CVA6Cfg[1092-:32] + 0))))) >= ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + (1 + (wbuffer_t_CVA6Cfg[1092-:32] + 0))))) ? ((wbuffer_t_CVA6Cfg[900-:32] + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + (wbuffer_t_CVA6Cfg[1092-:32] + 0))))) - ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + (1 + (wbuffer_t_CVA6Cfg[1092-:32] + 0)))))) + 1 : (((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + (1 + (wbuffer_t_CVA6Cfg[1092-:32] + 0))))) - (wbuffer_t_CVA6Cfg[900-:32] + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + (wbuffer_t_CVA6Cfg[1092-:32] + 0)))))) + 1)];
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:271:3
	assign wbuffer_be = (|wbuffer_hit_oh ? wbuffer_data_i[(wbuffer_hit_idx * ((((((((wbuffer_t_CVA6Cfg[996-:32] + (wbuffer_t_CVA6Cfg[1028-:32] - wbuffer_t_CVA6Cfg[9411 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9411 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9379 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9411 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9379 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9379 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9411 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)])) + wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)]) + wbuffer_t_CVA6Cfg[900-:32]) + (wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8)) + (wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8)) + (wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8)) + 1) + wbuffer_t_CVA6Cfg[1092-:32])) + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + (wbuffer_t_CVA6Cfg[1092-:32] + 0)))-:(((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + (wbuffer_t_CVA6Cfg[1092-:32] + 0))) >= ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + (1 + (wbuffer_t_CVA6Cfg[1092-:32] + 0))) ? (((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + (wbuffer_t_CVA6Cfg[1092-:32] + 0))) - ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + (1 + (wbuffer_t_CVA6Cfg[1092-:32] + 0)))) + 1 : (((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + (1 + (wbuffer_t_CVA6Cfg[1092-:32] + 0))) - ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + ((wbuffer_t_CVA6Cfg[9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))-:((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) >= (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) ? ((9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353))))))))) - (9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354)))))))))) + 1 : ((9509 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1354))))))))) - (9541 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + (32 + ((wbuffer_t_config_pkg_NrMaxRules * 64) + ((wbuffer_t_config_pkg_NrMaxRules * 64) + 1353)))))))))) + 1)] / 8) + (wbuffer_t_CVA6Cfg[1092-:32] + 0)))) + 1)] : {CVA6Cfg[17102-:32] / 8 {1'sb0}});
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:273:3
	generate
		if (CVA6Cfg[7625-:32] == 32'd0) begin : gen_axi_offset
			// Trace: core/cache_subsystem/wt_dcache_mem.sv:275:5
			assign wr_cl_off = (wr_cl_nc_i ? (CVA6Cfg[16712-:32] == CVA6Cfg[17102-:32] ? {CVA6Cfg[868-:32] - CVA6Cfg[16972-:32] {1'sb0}} : {{CVA6Cfg[868-:32] - AXI_OFFSET_WIDTH {1'b0}}, wr_cl_off_i[AXI_OFFSET_WIDTH - 1:CVA6Cfg[16972-:32]]}) : wr_cl_off_i[CVA6Cfg[868-:32] - 1:CVA6Cfg[16972-:32]]);
		end
		else begin : gen_piton_offset
			// Trace: core/cache_subsystem/wt_dcache_mem.sv:279:5
			assign wr_cl_off = wr_cl_off_i[CVA6Cfg[868-:32] - 1:3];
		end
	endgenerate
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:282:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: core/cache_subsystem/wt_dcache_mem.sv:283:5
		if (wr_cl_vld_i) begin
			// Trace: core/cache_subsystem/wt_dcache_mem.sv:284:7
			rdata = wr_cl_data_i[wr_cl_off * CVA6Cfg[17102-:32]+:CVA6Cfg[17102-:32]];
			// Trace: core/cache_subsystem/wt_dcache_mem.sv:285:7
			ruser = wr_cl_user_i[wr_cl_off * CVA6Cfg[900-:32]+:CVA6Cfg[900-:32]];
		end
		else begin
			// Trace: core/cache_subsystem/wt_dcache_mem.sv:287:7
			rdata = rdata_cl[rd_hit_idx * CVA6Cfg[17102-:32]+:CVA6Cfg[17102-:32]];
			// Trace: core/cache_subsystem/wt_dcache_mem.sv:288:7
			ruser = ruser_cl[rd_hit_idx * CVA6Cfg[900-:32]+:CVA6Cfg[900-:32]];
		end
	end
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:293:3
	genvar _gv_k_11;
	generate
		for (_gv_k_11 = 0; _gv_k_11 < (CVA6Cfg[17102-:32] / 8); _gv_k_11 = _gv_k_11 + 1) begin : gen_rd_data
			localparam k = _gv_k_11;
			// Trace: core/cache_subsystem/wt_dcache_mem.sv:294:5
			assign rd_data_o[8 * k+:8] = (wbuffer_be[k] ? wbuffer_rdata[8 * k+:8] : rdata[8 * k+:8]);
		end
	endgenerate
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:296:3
	genvar _gv_k_12;
	generate
		for (_gv_k_12 = 0; _gv_k_12 < (CVA6Cfg[900-:32] / 8); _gv_k_12 = _gv_k_12 + 1) begin : gen_rd_user
			localparam k = _gv_k_12;
			// Trace: core/cache_subsystem/wt_dcache_mem.sv:297:5
			assign rd_user_o[8 * k+:8] = (wbuffer_be[k] ? wbuffer_ruser[8 * k+:8] : ruser[8 * k+:8]);
		end
	endgenerate
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:304:3
	wire [CVA6Cfg[996-:32]:0] vld_tag_rdata [CVA6Cfg[1092-:32] - 1:0];
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:306:3
	genvar _gv_k_13;
	generate
		for (_gv_k_13 = 0; _gv_k_13 < DCACHE_NUM_BANKS; _gv_k_13 = _gv_k_13 + 1) begin : gen_data_banks
			localparam k = _gv_k_13;
			// Trace: core/cache_subsystem/wt_dcache_mem.sv:308:5
			sram_cache #(
				.USER_WIDTH(CVA6Cfg[1092-:32] * CVA6Cfg[900-:32]),
				.DATA_WIDTH(CVA6Cfg[1092-:32] * CVA6Cfg[17102-:32]),
				.USER_EN(CVA6Cfg[772-:32]),
				.BYTE_ACCESS(1),
				.TECHNO_CUT(CVA6Cfg[16875]),
				.NUM_WORDS(CVA6Cfg[836-:32])
			) i_data_sram(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.req_i(bank_req[k]),
				.we_i(bank_we[k]),
				.addr_i(bank_idx[k * DCACHE_CL_IDX_WIDTH+:DCACHE_CL_IDX_WIDTH]),
				.wuser_i(bank_wuser[CVA6Cfg[900-:32] * (k * CVA6Cfg[1092-:32])+:CVA6Cfg[900-:32] * CVA6Cfg[1092-:32]]),
				.wdata_i(bank_wdata[CVA6Cfg[17102-:32] * (k * CVA6Cfg[1092-:32])+:CVA6Cfg[17102-:32] * CVA6Cfg[1092-:32]]),
				.be_i(bank_be[(CVA6Cfg[17102-:32] / 8) * (k * CVA6Cfg[1092-:32])+:(CVA6Cfg[17102-:32] / 8) * CVA6Cfg[1092-:32]]),
				.ruser_o(bank_ruser[CVA6Cfg[900-:32] * (k * CVA6Cfg[1092-:32])+:CVA6Cfg[900-:32] * CVA6Cfg[1092-:32]]),
				.rdata_o(bank_rdata[CVA6Cfg[17102-:32] * (k * CVA6Cfg[1092-:32])+:CVA6Cfg[17102-:32] * CVA6Cfg[1092-:32]])
			);
		end
	endgenerate
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:329:3
	genvar _gv_i_70;
	generate
		for (_gv_i_70 = 0; _gv_i_70 < CVA6Cfg[1092-:32]; _gv_i_70 = _gv_i_70 + 1) begin : gen_tag_srams
			localparam i = _gv_i_70;
			// Trace: core/cache_subsystem/wt_dcache_mem.sv:331:5
			assign tag_rdata[i * CVA6Cfg[996-:32]+:CVA6Cfg[996-:32]] = vld_tag_rdata[i][CVA6Cfg[996-:32] - 1:0];
			// Trace: core/cache_subsystem/wt_dcache_mem.sv:332:5
			assign rd_vld_bits_o[i] = vld_tag_rdata[i][CVA6Cfg[996-:32]];
			// Trace: core/cache_subsystem/wt_dcache_mem.sv:335:5
			localparam sv2v_uu_i_tag_sram_USER_WIDTH = 1;
			// removed localparam type sv2v_uu_i_tag_sram_wuser_i
			localparam [0:0] sv2v_uu_i_tag_sram_ext_wuser_i_0 = 1'sb0;
			localparam sv2v_uu_i_tag_sram_DATA_WIDTH = CVA6Cfg[996-:32] + 1;
			// removed localparam type sv2v_uu_i_tag_sram_be_i
			localparam [((CVA6Cfg[996-:32] + 8) / 8) - 1:0] sv2v_uu_i_tag_sram_ext_be_i_1 = 1'sb1;
			sram_cache #(
				.DATA_WIDTH(CVA6Cfg[996-:32] + 1),
				.BYTE_ACCESS(0),
				.TECHNO_CUT(CVA6Cfg[16875]),
				.NUM_WORDS(CVA6Cfg[836-:32])
			) i_tag_sram(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.req_i(vld_req[i]),
				.we_i(vld_we),
				.addr_i(vld_addr),
				.wuser_i(sv2v_uu_i_tag_sram_ext_wuser_i_0),
				.wdata_i({vld_wdata[i], wr_cl_tag_i}),
				.be_i(sv2v_uu_i_tag_sram_ext_be_i_1),
				.ruser_o(),
				.rdata_o(vld_tag_rdata[i])
			);
		end
	endgenerate
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:355:3
	always @(posedge clk_i or negedge rst_ni) begin : p_regs
		// Trace: core/cache_subsystem/wt_dcache_mem.sv:356:5
		if (!rst_ni) begin
			// Trace: core/cache_subsystem/wt_dcache_mem.sv:357:7
			bank_idx_q <= 1'sb0;
			// Trace: core/cache_subsystem/wt_dcache_mem.sv:358:7
			bank_off_q <= 1'sb0;
			// Trace: core/cache_subsystem/wt_dcache_mem.sv:359:7
			vld_sel_q <= 1'sb0;
			// Trace: core/cache_subsystem/wt_dcache_mem.sv:360:7
			cmp_en_q <= 1'sb0;
		end
		else begin
			// Trace: core/cache_subsystem/wt_dcache_mem.sv:362:7
			bank_idx_q <= bank_idx_d;
			// Trace: core/cache_subsystem/wt_dcache_mem.sv:363:7
			bank_off_q <= bank_off_d;
			// Trace: core/cache_subsystem/wt_dcache_mem.sv:364:7
			vld_sel_q <= vld_sel_d;
			// Trace: core/cache_subsystem/wt_dcache_mem.sv:365:7
			cmp_en_q <= cmp_en_d;
		end
	end
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:375:3
	initial begin
		// Trace: core/cache_subsystem/wt_dcache_mem.sv:376:5
		begin : cach_line_width_axi
			
		end
	end
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:381:3
	initial begin
		// Trace: core/cache_subsystem/wt_dcache_mem.sv:382:5
		begin : axi_xlen
			
		end
	end
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:387:3
	initial begin
		// Trace: core/cache_subsystem/wt_dcache_mem.sv:388:5
		begin : cach_line_width_xlen
			
		end
	end
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:393:3
	// removed an assertion item
	// hit_hot1 : assert property (@(posedge clk_i) disable iff (!rst_ni)
	// 	(&vld_req |-> (!vld_we |=> $onehot0(rd_hit_oh_o)))
	// ) else begin
	// 	// Trace: core/cache_subsystem/wt_dcache_mem.sv:397:8
	// 	$fatal(1, "[l1 dcache] rd_hit_oh_o signal must be hot1");
	// end
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:399:3
	// removed an assertion item
	// word_write_hot1 : assert property (@(posedge clk_i) disable iff (!rst_ni)
	// 	(wr_ack_o |-> $onehot0(wr_req_i))
	// ) else begin
	// 	// Trace: core/cache_subsystem/wt_dcache_mem.sv:401:8
	// 	$fatal(1, "[l1 dcache] wr_req_i signal must be hot1");
	// end
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:403:3
	// removed an assertion item
	// wbuffer_hit_hot1 : assert property (@(posedge clk_i) disable iff (!rst_ni)
	// 	(&vld_req |-> (!vld_we |=> $onehot0(wbuffer_hit_oh)))
	// ) else begin
	// 	// Trace: core/cache_subsystem/wt_dcache_mem.sv:407:8
	// 	$fatal(1, "[l1 dcache] wbuffer_hit_oh signal must be hot1");
	// end
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:410:3
	reg [(CVA6Cfg[836-:32] * CVA6Cfg[1092-:32]) - 1:0] vld_mirror;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:411:3
	reg [((CVA6Cfg[836-:32] * CVA6Cfg[1092-:32]) * CVA6Cfg[996-:32]) - 1:0] tag_mirror;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:412:3
	wire [CVA6Cfg[1092-:32] - 1:0] tag_write_duplicate_test;
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:414:3
	function automatic [CVA6Cfg[1092-:32] - 1:0] sv2v_cast_B4195;
		input reg [CVA6Cfg[1092-:32] - 1:0] inp;
		sv2v_cast_B4195 = inp;
	endfunction
	function automatic [(CVA6Cfg[1092-:32] * CVA6Cfg[996-:32]) - 1:0] sv2v_cast_91A85;
		input reg [(CVA6Cfg[1092-:32] * CVA6Cfg[996-:32]) - 1:0] inp;
		sv2v_cast_91A85 = inp;
	endfunction
	always @(posedge clk_i or negedge rst_ni) begin : p_mirror
		// Trace: core/cache_subsystem/wt_dcache_mem.sv:415:5
		if (!rst_ni) begin
			// Trace: core/cache_subsystem/wt_dcache_mem.sv:416:7
			vld_mirror <= {CVA6Cfg[836-:32] {sv2v_cast_B4195(1'sb0)}};
			// Trace: core/cache_subsystem/wt_dcache_mem.sv:417:7
			tag_mirror <= {CVA6Cfg[836-:32] {sv2v_cast_91A85(1'sb0)}};
		end
		else
			// Trace: core/cache_subsystem/wt_dcache_mem.sv:419:7
			begin : sv2v_autoblock_2
				// Trace: core/cache_subsystem/wt_dcache_mem.sv:419:12
				reg signed [31:0] i;
				// Trace: core/cache_subsystem/wt_dcache_mem.sv:419:12
				for (i = 0; i < CVA6Cfg[1092-:32]; i = i + 1)
					begin
						// Trace: core/cache_subsystem/wt_dcache_mem.sv:420:9
						if (vld_req[i] & vld_we) begin
							// Trace: core/cache_subsystem/wt_dcache_mem.sv:421:11
							vld_mirror[(vld_addr * CVA6Cfg[1092-:32]) + i] <= vld_wdata[i];
							// Trace: core/cache_subsystem/wt_dcache_mem.sv:422:11
							tag_mirror[((vld_addr * CVA6Cfg[1092-:32]) + i) * CVA6Cfg[996-:32]+:CVA6Cfg[996-:32]] <= wr_cl_tag_i;
						end
					end
			end
	end
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:428:3
	genvar _gv_i_71;
	generate
		for (_gv_i_71 = 0; _gv_i_71 < CVA6Cfg[1092-:32]; _gv_i_71 = _gv_i_71 + 1) begin : gen_tag_dubl_test
			localparam i = _gv_i_71;
			// Trace: core/cache_subsystem/wt_dcache_mem.sv:429:5
			assign tag_write_duplicate_test[i] = ((tag_mirror[((vld_addr * CVA6Cfg[1092-:32]) + i) * CVA6Cfg[996-:32]+:CVA6Cfg[996-:32]] == wr_cl_tag_i) & vld_mirror[(vld_addr * CVA6Cfg[1092-:32]) + i]) & |vld_wdata;
		end
	endgenerate
	// Trace: core/cache_subsystem/wt_dcache_mem.sv:432:3
	// removed an assertion item
	// tag_write_duplicate : assert property (@(posedge clk_i) disable iff (!rst_ni)
	// 	(|vld_req |-> (vld_we |-> !(|tag_write_duplicate_test)))
	// ) else begin
	// 	// Trace: core/cache_subsystem/wt_dcache_mem.sv:435:8
	// 	$fatal(1, "[l1 dcache] cannot allocate a CL that is already present in the cache");
	// end
	initial _sv2v_0 = 0;
endmodule
