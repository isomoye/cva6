module cva6_rvfi_probes_5C276_3A398 (
	flush_i,
	issue_instr_ack_i,
	fetch_entry_valid_i,
	instruction_i,
	is_compressed_i,
	issue_pointer_i,
	commit_pointer_i,
	flush_unissued_instr_i,
	decoded_instr_valid_i,
	decoded_instr_ack_i,
	rs1_forwarding_i,
	rs2_forwarding_i,
	commit_instr_i,
	commit_drop_i,
	ex_commit_i,
	priv_lvl_i,
	lsu_ctrl_i,
	wbdata_i,
	commit_ack_i,
	mem_paddr_i,
	debug_mode_i,
	wdata_i,
	csr_i,
	rvfi_probes_o
);
	// removed localparam type exception_t_CVA6Cfg_type
	parameter [17102:0] exception_t_CVA6Cfg = 0;
	// removed localparam type lsu_ctrl_t_CVA6Cfg_type
	parameter [17102:0] lsu_ctrl_t_CVA6Cfg = 0;
	// removed localparam type scoreboard_entry_t_CVA6Cfg_type
	parameter [17102:0] scoreboard_entry_t_CVA6Cfg = 0;
	reg _sv2v_0;
	// removed import ariane_pkg::*;
	// Trace: core/cva6_rvfi_probes.sv:15:15
	localparam config_pkg_NrMaxRules = 16;
	// removed localparam type config_pkg_cache_type_t
	// removed localparam type config_pkg_noc_type_e
	// removed localparam type config_pkg_vm_mode_t
	// removed localparam type config_pkg_cva6_cfg_t
	localparam [17102:0] config_pkg_cva6_cfg_empty = 17103'd0;
	parameter [17102:0] CVA6Cfg = config_pkg_cva6_cfg_empty;
	// Trace: core/cva6_rvfi_probes.sv:16:20
	// removed localparam type exception_t
	// Trace: core/cva6_rvfi_probes.sv:17:20
	// removed localparam type scoreboard_entry_t
	// Trace: core/cva6_rvfi_probes.sv:18:20
	// removed localparam type lsu_ctrl_t
	// Trace: core/cva6_rvfi_probes.sv:19:20
	// removed localparam type rvfi_probes_instr_t
	// Trace: core/cva6_rvfi_probes.sv:20:20
	// removed localparam type rvfi_probes_csr_t
	// Trace: core/cva6_rvfi_probes.sv:21:20
	// removed localparam type rvfi_probes_t
	// Trace: core/cva6_rvfi_probes.sv:25:5
	input wire flush_i;
	// Trace: core/cva6_rvfi_probes.sv:26:5
	input wire [CVA6Cfg[16841-:32] - 1:0] issue_instr_ack_i;
	// Trace: core/cva6_rvfi_probes.sv:27:5
	input wire [CVA6Cfg[16841-:32] - 1:0] fetch_entry_valid_i;
	// Trace: core/cva6_rvfi_probes.sv:28:5
	input wire [(CVA6Cfg[16841-:32] * 32) - 1:0] instruction_i;
	// Trace: core/cva6_rvfi_probes.sv:29:5
	input wire [CVA6Cfg[16841-:32] - 1:0] is_compressed_i;
	// Trace: core/cva6_rvfi_probes.sv:31:5
	input wire [(CVA6Cfg[16841-:32] * CVA6Cfg[16503-:32]) - 1:0] issue_pointer_i;
	// Trace: core/cva6_rvfi_probes.sv:32:5
	input wire [(CVA6Cfg[16873-:32] * CVA6Cfg[16503-:32]) - 1:0] commit_pointer_i;
	// Trace: core/cva6_rvfi_probes.sv:34:5
	input wire flush_unissued_instr_i;
	// Trace: core/cva6_rvfi_probes.sv:35:5
	input wire [CVA6Cfg[16841-:32] - 1:0] decoded_instr_valid_i;
	// Trace: core/cva6_rvfi_probes.sv:36:5
	input wire [CVA6Cfg[16841-:32] - 1:0] decoded_instr_ack_i;
	// Trace: core/cva6_rvfi_probes.sv:38:5
	input wire [(CVA6Cfg[16841-:32] * CVA6Cfg[17070-:32]) - 1:0] rs1_forwarding_i;
	// Trace: core/cva6_rvfi_probes.sv:39:5
	input wire [(CVA6Cfg[16841-:32] * CVA6Cfg[17070-:32]) - 1:0] rs2_forwarding_i;
	// Trace: core/cva6_rvfi_probes.sv:41:5
	input wire [((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (CVA6Cfg[16873-:32] * (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5)) - 1 : (CVA6Cfg[16873-:32] * (1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 3)):((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 0 : ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)] commit_instr_i;
	// Trace: core/cva6_rvfi_probes.sv:42:5
	input wire [CVA6Cfg[16873-:32] - 1:0] commit_drop_i;
	// Trace: core/cva6_rvfi_probes.sv:43:5
	input wire [((exception_t_CVA6Cfg[17102-:32] + exception_t_CVA6Cfg[17102-:32]) + exception_t_CVA6Cfg[17006-:32]) + 33:0] ex_commit_i;
	// Trace: core/cva6_rvfi_probes.sv:44:5
	// removed localparam type riscv_priv_lvl_t
	input wire [1:0] priv_lvl_i;
	// Trace: core/cva6_rvfi_probes.sv:46:5
	input wire [((((((1 + lsu_ctrl_t_CVA6Cfg[17070-:32]) + 36) + lsu_ctrl_t_CVA6Cfg[17102-:32]) + (lsu_ctrl_t_CVA6Cfg[17102-:32] / 8)) + 12) + lsu_ctrl_t_CVA6Cfg[16503-:32]) - 1:0] lsu_ctrl_i;
	// Trace: core/cva6_rvfi_probes.sv:47:5
	input wire [(CVA6Cfg[16401-:32] * CVA6Cfg[17102-:32]) - 1:0] wbdata_i;
	// Trace: core/cva6_rvfi_probes.sv:48:5
	input wire [CVA6Cfg[16873-:32] - 1:0] commit_ack_i;
	// Trace: core/cva6_rvfi_probes.sv:49:5
	input wire [CVA6Cfg[17038-:32] - 1:0] mem_paddr_i;
	// Trace: core/cva6_rvfi_probes.sv:50:5
	input wire debug_mode_i;
	// Trace: core/cva6_rvfi_probes.sv:51:5
	input wire [(CVA6Cfg[16873-:32] * CVA6Cfg[17102-:32]) - 1:0] wdata_i;
	// Trace: core/cva6_rvfi_probes.sv:53:5
	input wire csr_i;
	// Trace: core/cva6_rvfi_probes.sv:55:5
	output reg [1:0] rvfi_probes_o;
	// Trace: core/cva6_rvfi_probes.sv:59:3
	reg csr;
	// Trace: core/cva6_rvfi_probes.sv:60:3
	reg instr;
	// Trace: core/cva6_rvfi_probes.sv:62:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: core/cva6_rvfi_probes.sv:63:5
		csr = 1'sb0;
		// Trace: core/cva6_rvfi_probes.sv:64:5
		instr = 1'sb0;
		// Trace: core/cva6_rvfi_probes.sv:66:5
		instr.flush = flush_i;
		// Trace: core/cva6_rvfi_probes.sv:67:5
		instr.issue_instr_ack = issue_instr_ack_i;
		// Trace: core/cva6_rvfi_probes.sv:68:5
		instr.fetch_entry_valid = fetch_entry_valid_i;
		// Trace: core/cva6_rvfi_probes.sv:69:5
		instr.instruction = instruction_i;
		// Trace: core/cva6_rvfi_probes.sv:70:5
		instr.is_compressed = is_compressed_i;
		// Trace: core/cva6_rvfi_probes.sv:72:5
		instr.issue_pointer = issue_pointer_i;
		// Trace: core/cva6_rvfi_probes.sv:74:5
		instr.flush_unissued_instr = flush_unissued_instr_i;
		// Trace: core/cva6_rvfi_probes.sv:75:5
		instr.decoded_instr_valid = decoded_instr_valid_i;
		// Trace: core/cva6_rvfi_probes.sv:76:5
		instr.decoded_instr_ack = decoded_instr_ack_i;
		// Trace: core/cva6_rvfi_probes.sv:78:5
		instr.rs1_forwarding = rs1_forwarding_i;
		// Trace: core/cva6_rvfi_probes.sv:79:5
		instr.rs2_forwarding = rs2_forwarding_i;
		// Trace: core/cva6_rvfi_probes.sv:81:5
		instr.ex_commit_cause = ex_commit_i[exception_t_CVA6Cfg[17102-:32] + (exception_t_CVA6Cfg[17102-:32] + (exception_t_CVA6Cfg[17006-:32] + 33))-:((exception_t_CVA6Cfg[17102-:32] + (exception_t_CVA6Cfg[17102-:32] + (exception_t_CVA6Cfg[17006-:32] + 33))) >= (exception_t_CVA6Cfg[17102-:32] + (exception_t_CVA6Cfg[17006-:32] + 34)) ? ((exception_t_CVA6Cfg[17102-:32] + (exception_t_CVA6Cfg[17102-:32] + (exception_t_CVA6Cfg[17006-:32] + 33))) - (exception_t_CVA6Cfg[17102-:32] + (exception_t_CVA6Cfg[17006-:32] + 34))) + 1 : ((exception_t_CVA6Cfg[17102-:32] + (exception_t_CVA6Cfg[17006-:32] + 34)) - (exception_t_CVA6Cfg[17102-:32] + (exception_t_CVA6Cfg[17102-:32] + (exception_t_CVA6Cfg[17006-:32] + 33)))) + 1)];
		// Trace: core/cva6_rvfi_probes.sv:82:5
		instr.ex_commit_valid = ex_commit_i[0];
		// Trace: core/cva6_rvfi_probes.sv:84:5
		instr.priv_lvl = priv_lvl_i;
		// Trace: core/cva6_rvfi_probes.sv:86:5
		instr.lsu_ctrl_vaddr = lsu_ctrl_i[lsu_ctrl_t_CVA6Cfg[17070-:32] + (36 + (lsu_ctrl_t_CVA6Cfg[17102-:32] + ((lsu_ctrl_t_CVA6Cfg[17102-:32] / 8) + (lsu_ctrl_t_CVA6Cfg[16503-:32] + 11))))-:((lsu_ctrl_t_CVA6Cfg[17070-:32] + (36 + (lsu_ctrl_t_CVA6Cfg[17102-:32] + ((lsu_ctrl_t_CVA6Cfg[17102-:32] / 8) + (lsu_ctrl_t_CVA6Cfg[16503-:32] + 11))))) >= (36 + (lsu_ctrl_t_CVA6Cfg[17102-:32] + ((lsu_ctrl_t_CVA6Cfg[17102-:32] / 8) + (12 + (lsu_ctrl_t_CVA6Cfg[16503-:32] + 0))))) ? ((lsu_ctrl_t_CVA6Cfg[17070-:32] + (36 + (lsu_ctrl_t_CVA6Cfg[17102-:32] + ((lsu_ctrl_t_CVA6Cfg[17102-:32] / 8) + (lsu_ctrl_t_CVA6Cfg[16503-:32] + 11))))) - (36 + (lsu_ctrl_t_CVA6Cfg[17102-:32] + ((lsu_ctrl_t_CVA6Cfg[17102-:32] / 8) + (12 + (lsu_ctrl_t_CVA6Cfg[16503-:32] + 0)))))) + 1 : ((36 + (lsu_ctrl_t_CVA6Cfg[17102-:32] + ((lsu_ctrl_t_CVA6Cfg[17102-:32] / 8) + (12 + (lsu_ctrl_t_CVA6Cfg[16503-:32] + 0))))) - (lsu_ctrl_t_CVA6Cfg[17070-:32] + (36 + (lsu_ctrl_t_CVA6Cfg[17102-:32] + ((lsu_ctrl_t_CVA6Cfg[17102-:32] / 8) + (lsu_ctrl_t_CVA6Cfg[16503-:32] + 11)))))) + 1)];
		// Trace: core/cva6_rvfi_probes.sv:87:5
		instr.lsu_ctrl_fu = lsu_ctrl_i[lsu_ctrl_t_CVA6Cfg[16503-:32] + 11-:((lsu_ctrl_t_CVA6Cfg[16503-:32] + 11) >= (8 + (lsu_ctrl_t_CVA6Cfg[16503-:32] + 0)) ? ((lsu_ctrl_t_CVA6Cfg[16503-:32] + 11) - (8 + (lsu_ctrl_t_CVA6Cfg[16503-:32] + 0))) + 1 : ((8 + (lsu_ctrl_t_CVA6Cfg[16503-:32] + 0)) - (lsu_ctrl_t_CVA6Cfg[16503-:32] + 11)) + 1)];
		// Trace: core/cva6_rvfi_probes.sv:88:5
		instr.lsu_ctrl_be = lsu_ctrl_i[(lsu_ctrl_t_CVA6Cfg[17102-:32] / 8) + (lsu_ctrl_t_CVA6Cfg[16503-:32] + 11)-:(((lsu_ctrl_t_CVA6Cfg[17102-:32] / 8) + (lsu_ctrl_t_CVA6Cfg[16503-:32] + 11)) >= (12 + (lsu_ctrl_t_CVA6Cfg[16503-:32] + 0)) ? (((lsu_ctrl_t_CVA6Cfg[17102-:32] / 8) + (lsu_ctrl_t_CVA6Cfg[16503-:32] + 11)) - (12 + (lsu_ctrl_t_CVA6Cfg[16503-:32] + 0))) + 1 : ((12 + (lsu_ctrl_t_CVA6Cfg[16503-:32] + 0)) - ((lsu_ctrl_t_CVA6Cfg[17102-:32] / 8) + (lsu_ctrl_t_CVA6Cfg[16503-:32] + 11))) + 1)];
		// Trace: core/cva6_rvfi_probes.sv:89:5
		instr.lsu_ctrl_trans_id = lsu_ctrl_i[lsu_ctrl_t_CVA6Cfg[16503-:32] - 1-:lsu_ctrl_t_CVA6Cfg[16503-:32]];
		// Trace: core/cva6_rvfi_probes.sv:91:5
		instr.wbdata = wbdata_i;
		// Trace: core/cva6_rvfi_probes.sv:92:5
		instr.mem_paddr = mem_paddr_i;
		// Trace: core/cva6_rvfi_probes.sv:93:5
		instr.debug_mode = debug_mode_i;
		// Trace: core/cva6_rvfi_probes.sv:95:5
		instr.commit_pointer = commit_pointer_i;
		// Trace: core/cva6_rvfi_probes.sv:97:5
		begin : sv2v_autoblock_1
			// Trace: core/cva6_rvfi_probes.sv:97:10
			reg signed [31:0] i;
			// Trace: core/cva6_rvfi_probes.sv:97:10
			for (i = 0; i < CVA6Cfg[16873-:32]; i = i + 1)
				begin
					// Trace: core/cva6_rvfi_probes.sv:98:7
					instr.commit_instr_pc[i] = commit_instr_i[((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? scoreboard_entry_t_CVA6Cfg[17070-:32] + (scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (scoreboard_entry_t_CVA6Cfg[17070-:32] + (scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))))) : (((i * ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? scoreboard_entry_t_CVA6Cfg[17070-:32] + (scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (scoreboard_entry_t_CVA6Cfg[17070-:32] + (scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))))) + ((scoreboard_entry_t_CVA6Cfg[17070-:32] + (scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) >= (scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) ? ((scoreboard_entry_t_CVA6Cfg[17070-:32] + (scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) - (scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))))) + 1 : ((scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) - (scoreboard_entry_t_CVA6Cfg[17070-:32] + (scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))))) + 1)) - 1)-:((scoreboard_entry_t_CVA6Cfg[17070-:32] + (scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) >= (scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) ? ((scoreboard_entry_t_CVA6Cfg[17070-:32] + (scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) - (scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))))) + 1 : ((scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) - (scoreboard_entry_t_CVA6Cfg[17070-:32] + (scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))))) + 1)];
					// Trace: core/cva6_rvfi_probes.sv:99:7
					instr.commit_instr_op[i] = commit_instr_i[((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((i * ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((23 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((23 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)];
					// Trace: core/cva6_rvfi_probes.sv:100:7
					instr.commit_instr_rs1[i] = commit_instr_i[((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 15 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (15 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((i * ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 15 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (15 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((15 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (10 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((15 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (10 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((10 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (15 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((15 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (10 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((15 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (10 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((10 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (15 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)];
					// Trace: core/cva6_rvfi_probes.sv:101:7
					instr.commit_instr_rs2[i] = commit_instr_i[((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 10 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (10 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((i * ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 10 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (10 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((10 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (5 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((10 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (5 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((5 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (10 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((10 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (5 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((10 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (5 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((5 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (10 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)];
					// Trace: core/cva6_rvfi_probes.sv:102:7
					instr.commit_instr_rd[i] = commit_instr_i[((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 5 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (5 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((i * ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 5 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (5 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((5 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) ? ((5 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) + 1 : ((scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) - (5 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((5 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) ? ((5 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) + 1 : ((scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) - (5 + (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)];
					// Trace: core/cva6_rvfi_probes.sv:103:7
					instr.commit_instr_result[i] = commit_instr_i[((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))) : (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) : (((i * ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))) : (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + ((scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) >= (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))) ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) + 1 : ((4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))) - (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + 1)) - 1)-:((scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) >= (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))) ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) + 1 : ((4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))) - (scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + 1)];
					// Trace: core/cva6_rvfi_probes.sv:104:7
					instr.commit_instr_valid[i] = commit_instr_i[(i * ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) : (((((((scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (4 + (((((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))];
				end
		end
		// Trace: core/cva6_rvfi_probes.sv:107:5
		instr.commit_drop = commit_drop_i;
		// Trace: core/cva6_rvfi_probes.sv:108:5
		instr.commit_ack = commit_ack_i;
		// Trace: core/cva6_rvfi_probes.sv:109:5
		instr.wdata = wdata_i;
		// Trace: core/cva6_rvfi_probes.sv:111:5
		csr = csr_i;
	end
	// Trace: core/cva6_rvfi_probes.sv:116:3
	always @(*) begin
		if (_sv2v_0)
			;
		// Trace: core/cva6_rvfi_probes.sv:117:5
		rvfi_probes_o = 1'sb0;
		// Trace: core/cva6_rvfi_probes.sv:119:5
		// Trace: core/cva6_rvfi_probes.sv:120:7
		rvfi_probes_o[0] = instr;
		// Trace: core/cva6_rvfi_probes.sv:124:7
		rvfi_probes_o[1] = csr;
	end
	initial _sv2v_0 = 0;
endmodule
