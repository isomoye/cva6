module cva6_hpdcache_if_adapter_D71A0_F1924 (
	clk_i,
	rst_ni,
	hpdcache_req_sid_i,
	cva6_req_i,
	cva6_req_o,
	cva6_amo_req_i,
	cva6_amo_resp_o,
	hpdcache_req_valid_o,
	hpdcache_req_ready_i,
	hpdcache_req_o,
	hpdcache_req_abort_o,
	hpdcache_req_tag_o,
	hpdcache_req_pma_o,
	hpdcache_rsp_valid_i,
	hpdcache_rsp_i
);
	// removed localparam type dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg_type
	parameter [17102:0] dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg = 0;
	// removed localparam type dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg_type
	parameter [17102:0] dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg = 0;
	// removed localparam type hpdcache_req_offset_t_hpdcache_req_offset_t_HPDcacheCfg_type
	parameter [1349:0] hpdcache_req_offset_t_hpdcache_req_offset_t_HPDcacheCfg = 0;
	// removed localparam type hpdcache_req_sid_t_hpdcache_req_sid_t_HPDcacheCfg_type
	parameter [1349:0] hpdcache_req_sid_t_hpdcache_req_sid_t_HPDcacheCfg = 0;
	// removed localparam type hpdcache_req_t_hpdcache_req_t_HPDcacheCfg_type
	parameter [1349:0] hpdcache_req_t_hpdcache_req_t_HPDcacheCfg = 0;
	// removed localparam type hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg_type
	parameter [1349:0] hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg = 0;
	// removed localparam type hpdcache_tag_t_hpdcache_tag_t_HPDcacheCfg_type
	parameter [1349:0] hpdcache_tag_t_hpdcache_tag_t_HPDcacheCfg = 0;
	reg _sv2v_0;
	// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:16:15
	localparam config_pkg_NrMaxRules = 16;
	// removed localparam type config_pkg_cache_type_t
	// removed localparam type config_pkg_noc_type_e
	// removed localparam type config_pkg_vm_mode_t
	// removed localparam type config_pkg_cva6_cfg_t
	localparam [17102:0] config_pkg_cva6_cfg_empty = 17103'd0;
	parameter [17102:0] CVA6Cfg = config_pkg_cva6_cfg_empty;
	// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:17:15
	// removed localparam type hpdcache_pkg_hpdcache_victim_sel_policy_t
	// removed localparam type hpdcache_pkg_hpdcache_user_cfg_t
	// removed localparam type hpdcache_pkg_hpdcache_cfg_t
	parameter [1349:0] HPDcacheCfg = 1'sb0;
	// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:18:20
	// removed localparam type hpdcache_tag_t
	// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:19:20
	// removed localparam type hpdcache_req_offset_t
	// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:20:20
	// removed localparam type hpdcache_req_sid_t
	// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:21:20
	// removed localparam type hpdcache_req_t
	// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:22:20
	// removed localparam type hpdcache_rsp_t
	// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:23:20
	// removed localparam type dcache_req_i_t
	// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:24:20
	// removed localparam type dcache_req_o_t
	// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:25:15
	parameter [0:0] is_load_port = 1'b1;
	// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:33:5
	input wire clk_i;
	// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:34:5
	input wire rst_ni;
	// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:37:5
	input wire [hpdcache_req_sid_t_hpdcache_req_sid_t_HPDcacheCfg[1093-:32] - 1:0] hpdcache_req_sid_i;
	// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:40:5
	input wire [(((((((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1028-:32] + dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[996-:32]) + dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32]) + dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32]) + 2) + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8)) + 2) + dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32]) + 1:0] cva6_req_i;
	// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:41:5
	output wire [(((2 + dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[1124-:32]) + dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[17102-:32]) + dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[900-:32]) - 1:0] cva6_req_o;
	// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:42:5
	// removed localparam type ariane_pkg_amo_t
	// removed localparam type ariane_pkg_amo_req_t
	input wire [134:0] cva6_amo_req_i;
	// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:43:5
	// removed localparam type ariane_pkg_amo_resp_t
	output wire [64:0] cva6_amo_resp_o;
	// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:46:5
	output wire hpdcache_req_valid_o;
	// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:47:5
	input wire hpdcache_req_ready_i;
	// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:48:5
	output wire [((((((((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32])) + 4) + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8))) + 3) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32]) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32]) + 2) + hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32]) + 1:0] hpdcache_req_o;
	// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:49:5
	output wire hpdcache_req_abort_o;
	// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:50:5
	output wire [hpdcache_tag_t_hpdcache_tag_t_HPDcacheCfg[351-:32] - 1:0] hpdcache_req_tag_o;
	// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:51:5
	// removed localparam type hpdcache_pkg_hpdcache_pma_t
	output wire [1:0] hpdcache_req_pma_o;
	// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:54:5
	input wire hpdcache_rsp_valid_i;
	// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:55:5
	input wire [(((hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1157-:32] * hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1285-:32]) + hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32]) + hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32]) + 1:0] hpdcache_rsp_i;
	// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:61:3
	wire forward_store;
	wire forward_amo;
	// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:62:3
	wire hpdcache_req_is_uncacheable;
	// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:67:3
	function automatic [64:0] sv2v_cast_65;
		input reg [64:0] inp;
		sv2v_cast_65 = inp;
	endfunction
	function automatic config_pkg_range_check;
		// Trace: core/include/config_pkg.sv:375:40
		input reg [63:0] base;
		// Trace: core/include/config_pkg.sv:375:59
		input reg [63:0] len;
		// Trace: core/include/config_pkg.sv:375:77
		input reg [63:0] address;
		// Trace: core/include/config_pkg.sv:378:5
		config_pkg_range_check = (address >= base) && ({1'b0, address} < (sv2v_cast_65(base) + len));
	endfunction
	function automatic config_pkg_is_inside_cacheable_regions;
		// Trace: core/include/config_pkg.sv:405:56
		input reg [17102:0] Cfg;
		// Trace: core/include/config_pkg.sv:405:72
		input reg [63:0] address;
		// Trace: core/include/config_pkg.sv:406:5
		reg [15:0] pass;
		begin
			// Trace: core/include/config_pkg.sv:407:5
			pass = 1'sb0;
			// Trace: core/include/config_pkg.sv:408:5
			begin : sv2v_autoblock_1
				// Trace: core/include/config_pkg.sv:408:10
				reg [31:0] k;
				// Trace: core/include/config_pkg.sv:408:10
				for (k = 0; k < Cfg[3433-:32]; k = k + 1)
					begin
						// Trace: core/include/config_pkg.sv:409:7
						pass[k] = config_pkg_range_check(Cfg[2378 + (k * 64)+:64], Cfg[1354 + (k * 64)+:64], address);
					end
			end
			config_pkg_is_inside_cacheable_regions = |pass;
		end
	endfunction
	// removed localparam type hpdcache_pkg_hpdcache_req_op_t
	generate
		if (is_load_port == 1'b1) begin : load_port_gen
			// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:71:7
			assign hpdcache_req_is_uncacheable = !config_pkg_is_inside_cacheable_regions(CVA6Cfg, {{64 - CVA6Cfg[996-:32] {1'b0}}, cva6_req_i[dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[996-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1))))))-:((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[996-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1))))))) >= (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2)))))) ? ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[996-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1))))))) - (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2))))))) + 1 : ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2)))))) - (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[996-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1)))))))) + 1)], {CVA6Cfg[1028-:32] {1'b0}}});
			// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:81:7
			assign hpdcache_req_valid_o = cva6_req_i[2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1)))];
			assign hpdcache_req_o[hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))-:((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))) >= ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))))) ? ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))) - ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))))) + 1 : (((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))))) - (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))))) + 1)] = cva6_req_i[dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1028-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[996-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1)))))))-:((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1028-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[996-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1)))))))) >= (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[996-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2))))))) ? ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1028-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[996-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1)))))))) - (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[996-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2)))))))) + 1 : ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[996-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2))))))) - (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1028-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[996-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1))))))))) + 1)];
			assign hpdcache_req_o[(hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))-:(((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) >= (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) ? (((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) - (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))))) + 1 : ((4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) - ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))) + 1)] = 1'sb0;
			assign hpdcache_req_o[4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))-:((4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) >= ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) ? ((4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) - ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) + 1 : (((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) - (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) + 1)] = 4'h0;
			assign hpdcache_req_o[(hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))-:(((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) >= (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))) ? (((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) - (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) + 1 : ((3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))) - ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) + 1)] = cva6_req_i[(dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1))-:(((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1))) >= (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2)) ? (((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1))) - (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2))) + 1 : ((2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2)) - ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1)))) + 1)];
			assign hpdcache_req_o[3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))-:((3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) >= (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) ? ((3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) - (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))) + 1 : ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) - (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) + 1)] = cva6_req_i[2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1)-:((2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1)) >= (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2) ? ((2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1)) - (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2)) + 1 : ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2) - (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1))) + 1)];
			assign hpdcache_req_o[hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))-:((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))) >= (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))) ? ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))) - (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) + 1 : ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))) - (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) + 1)] = hpdcache_req_sid_i;
			assign hpdcache_req_o[hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))-:((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))) >= (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)) ? ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))) - (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))) + 1 : ((2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)) - (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))) + 1)] = cva6_req_i[dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1-:((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1) >= 2 ? dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 0 : 3 - (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1))];
			assign hpdcache_req_o[2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)] = 1'b1;
			assign hpdcache_req_o[1 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)] = 1'b0;
			assign hpdcache_req_o[hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1-:((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1) >= 2 ? hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 0 : 3 - (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))] = 1'sb0;
			assign hpdcache_req_o[1-:2] = 1'sb0;
			// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:94:7
			assign hpdcache_req_abort_o = cva6_req_i[1];
			assign hpdcache_req_tag_o = cva6_req_i[dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[996-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1))))))-:((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[996-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1))))))) >= (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2)))))) ? ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[996-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1))))))) - (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2))))))) + 1 : ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2)))))) - (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[996-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1)))))))) + 1)];
			assign hpdcache_req_pma_o[1] = hpdcache_req_is_uncacheable;
			assign hpdcache_req_pma_o[0] = 1'b0;
			// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:100:7
			assign cva6_req_o[1 + (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[1124-:32] + (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[17102-:32] + (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[900-:32] - 1)))] = hpdcache_rsp_valid_i;
			assign cva6_req_o[dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[17102-:32] + (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[900-:32] - 1)-:((dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[17102-:32] + (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[900-:32] - 1)) >= (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[900-:32] + 0) ? ((dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[17102-:32] + (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[900-:32] - 1)) - (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[900-:32] + 0)) + 1 : ((dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[900-:32] + 0) - (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[17102-:32] + (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[900-:32] - 1))) + 1)] = hpdcache_rsp_i[(hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1157-:32] * hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1285-:32]) + (hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32] + (hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1))-:(((hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1157-:32] * hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1285-:32]) + (hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32] + (hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1))) >= (hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32] + (hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 2)) ? (((hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1157-:32] * hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1285-:32]) + (hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32] + (hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1))) - (hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32] + (hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 2))) + 1 : ((hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32] + (hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 2)) - ((hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1157-:32] * hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1285-:32]) + (hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32] + (hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1)))) + 1)];
			assign cva6_req_o[dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[1124-:32] + (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[17102-:32] + (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[900-:32] - 1))-:((dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[1124-:32] + (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[17102-:32] + (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[900-:32] - 1))) >= (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[17102-:32] + (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[900-:32] + 0)) ? ((dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[1124-:32] + (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[17102-:32] + (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[900-:32] - 1))) - (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[17102-:32] + (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[900-:32] + 0))) + 1 : ((dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[17102-:32] + (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[900-:32] + 0)) - (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[1124-:32] + (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[17102-:32] + (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[900-:32] - 1)))) + 1)] = hpdcache_rsp_i[hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1-:((hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1) >= 2 ? hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 0 : 3 - (hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1))];
			assign cva6_req_o[2 + (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[1124-:32] + (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[17102-:32] + (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[900-:32] - 1)))] = hpdcache_req_ready_i;
		end
		else begin : store_amo_gen
			// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:109:7
			reg [63:0] amo_addr;
			// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:110:7
			reg [hpdcache_req_offset_t_hpdcache_req_offset_t_HPDcacheCfg[287-:32] - 1:0] amo_addr_offset;
			// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:111:7
			reg [hpdcache_tag_t_hpdcache_tag_t_HPDcacheCfg[351-:32] - 1:0] amo_tag;
			// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:112:7
			wire amo_is_word;
			wire amo_is_word_hi;
			// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:113:7
			wire [63:0] amo_data;
			// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:114:7
			wire [7:0] amo_data_be;
			// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:115:7
			reg [3:0] amo_op;
			// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:116:7
			wire [31:0] amo_resp_word;
			// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:117:7
			reg amo_pending_q;
			// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:121:7
			always @(*) begin : amo_op_comb
				if (_sv2v_0)
					;
				// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:122:9
				amo_addr = cva6_amo_req_i[127-:64];
				// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:123:9
				amo_addr_offset = amo_addr[0+:HPDcacheCfg[287-:32]];
				// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:124:9
				amo_tag = amo_addr[HPDcacheCfg[287-:32]+:HPDcacheCfg[351-:32]];
				// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:125:9
				(* full_case, parallel_case *)
				case (cva6_amo_req_i[133-:4])
					4'b0001:
						// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:126:33
						amo_op = 4'h4;
					4'b0010:
						// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:127:33
						amo_op = 4'h5;
					4'b0011:
						// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:128:33
						amo_op = 4'h6;
					4'b0100:
						// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:129:33
						amo_op = 4'h7;
					4'b0101:
						// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:130:33
						amo_op = 4'h8;
					4'b0110:
						// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:131:33
						amo_op = 4'h9;
					4'b0111:
						// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:132:33
						amo_op = 4'ha;
					4'b1000:
						// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:133:33
						amo_op = 4'hb;
					4'b1001:
						// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:134:33
						amo_op = 4'hc;
					4'b1010:
						// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:135:33
						amo_op = 4'hd;
					4'b1011:
						// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:136:33
						amo_op = 4'he;
					default:
						// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:137:33
						amo_op = 4'h0;
				endcase
			end
			// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:144:7
			assign hpdcache_req_is_uncacheable = !config_pkg_is_inside_cacheable_regions(CVA6Cfg, {{64 - CVA6Cfg[996-:32] {1'b0}}, hpdcache_req_o[hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1-:((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1) >= 2 ? hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 0 : 3 - (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))], {CVA6Cfg[1028-:32] {1'b0}}});
			// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:153:7
			assign amo_is_word = cva6_amo_req_i[129-:2] == 2'b10;
			// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:154:7
			assign amo_is_word_hi = cva6_amo_req_i[66];
			if (CVA6Cfg[17102-:32] == 64) begin : amo_data_64_gen
				// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:156:9
				assign amo_data = (amo_is_word ? {2 {cva6_amo_req_i[0+:32]}} : cva6_amo_req_i[63-:64]);
				// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:157:9
				assign amo_data_be = (amo_is_word_hi ? 8'hf0 : (amo_is_word ? 8'h0f : 8'hff));
			end
			else begin : amo_data_32_gen
				// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:159:9
				assign amo_data = {32'b00000000000000000000000000000000, cva6_amo_req_i[63-:64]};
				// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:160:9
				assign amo_data_be = 8'h0f;
			end
			// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:163:7
			assign forward_store = cva6_req_i[2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1)))];
			// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:164:7
			assign forward_amo = cva6_amo_req_i[134];
			// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:166:7
			assign hpdcache_req_valid_o = forward_store | (forward_amo & ~amo_pending_q);
			// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:167:7
			assign hpdcache_req_o[hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))-:((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))) >= ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))))) ? ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))) - ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))))) + 1 : (((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))))) - (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[287-:32] + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))))) + 1)] = (forward_amo ? amo_addr_offset : cva6_req_i[dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1028-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[996-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1)))))))-:((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1028-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[996-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1)))))))) >= (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[996-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2))))))) ? ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1028-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[996-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1)))))))) - (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[996-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2)))))))) + 1 : ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[996-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2))))))) - (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1028-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[996-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1))))))))) + 1)]);
			// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:168:7
			assign hpdcache_req_o[(hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))-:(((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) >= (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) ? (((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) - (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))))) + 1 : ((4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) - ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32]) + (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))))) + 1)] = (forward_amo ? amo_data : cva6_req_i[dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1)))))-:((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1)))))) >= (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2))))) ? ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1)))))) - (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2)))))) + 1 : ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2))))) - (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1))))))) + 1)]);
			// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:169:7
			assign hpdcache_req_o[4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))-:((4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) >= ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) ? ((4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) - ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))))) + 1 : (((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) - (4 + ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))))) + 1)] = (forward_amo ? amo_op : 4'h1);
			// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:170:7
			assign hpdcache_req_o[(hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))-:(((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) >= (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))) ? (((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) - (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))))) + 1 : ((3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))) - ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1157-:32] * (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1285-:32] / 8)) + (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))))) + 1)] = (forward_amo ? amo_data_be : cva6_req_i[(dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1))-:(((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1))) >= (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2)) ? (((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1))) - (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2))) + 1 : ((2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2)) - ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1)))) + 1)]);
			// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:171:7
			assign hpdcache_req_o[3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))-:((3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) >= (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) ? ((3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) - (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))))) + 1 : ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) - (3 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))))) + 1)] = (forward_amo ? cva6_amo_req_i[129-:2] : cva6_req_i[2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1)-:((2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1)) >= (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2) ? ((2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1)) - (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2)) + 1 : ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2) - (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1))) + 1)]);
			// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:172:7
			assign hpdcache_req_o[hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))-:((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))) >= (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))) ? ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))) - (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)))) + 1 : ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))) - (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1093-:32] + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))))) + 1)] = hpdcache_req_sid_i;
			// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:173:7
			assign hpdcache_req_o[hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))-:((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))) >= (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)) ? ((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))) - (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2))) + 1 : ((2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 2)) - (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] + (2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)))) + 1)] = (forward_amo ? {hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] {1'sb1}} : {hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[1125-:32] {1'sb0}});
			// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:174:7
			assign hpdcache_req_o[2 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)] = forward_amo;
			// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:175:7
			assign hpdcache_req_o[1 + (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1)] = 1'b1;
			// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:176:7
			assign hpdcache_req_o[hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1-:((hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1) >= 2 ? hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 0 : 3 - (hpdcache_req_t_hpdcache_req_t_HPDcacheCfg[351-:32] + 1))] = (forward_amo ? amo_tag : cva6_req_i[dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[996-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1))))))-:((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[996-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1))))))) >= (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2)))))) ? ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[996-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1))))))) - (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2))))))) + 1 : ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2)))))) - (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[996-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1)))))))) + 1)]);
			// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:177:7
			assign hpdcache_req_o[1] = hpdcache_req_is_uncacheable;
			// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:178:7
			assign hpdcache_req_o[0] = 1'b0;
			// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:179:7
			assign hpdcache_req_abort_o = 1'b0;
			// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:180:7
			assign hpdcache_req_tag_o = 1'sb0;
			// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:181:7
			assign hpdcache_req_pma_o = 1'sb0;
			if (CVA6Cfg[17102-:32] == 64) begin : amo_resp_64_gen
				// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:187:9
				assign amo_resp_word = (amo_is_word_hi ? hpdcache_rsp_i[((hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1157-:32] * hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1285-:32]) + (hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32] + (hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1))) - ((hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1157-:32] * hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1285-:32]) - 33)+:32] : hpdcache_rsp_i[((hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1157-:32] * hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1285-:32]) + (hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32] + (hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1))) - ((hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1157-:32] * hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1285-:32]) - 1)+:32]);
			end
			else begin : amo_resp_32_gen
				// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:191:9
				assign amo_resp_word = hpdcache_rsp_i[((hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1157-:32] * hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1285-:32]) + (hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32] + (hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1))) - ((hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1157-:32] * hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1285-:32]) - 1)+:hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1285-:32]];
			end
			// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:194:7
			assign cva6_req_o[1 + (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[1124-:32] + (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[17102-:32] + (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[900-:32] - 1)))] = hpdcache_rsp_valid_i && (hpdcache_rsp_i[hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1-:((hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1) >= 2 ? hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 0 : 3 - (hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1))] != {hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] {1'sb1}});
			// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:195:7
			assign cva6_req_o[dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[17102-:32] + (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[900-:32] - 1)-:((dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[17102-:32] + (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[900-:32] - 1)) >= (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[900-:32] + 0) ? ((dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[17102-:32] + (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[900-:32] - 1)) - (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[900-:32] + 0)) + 1 : ((dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[900-:32] + 0) - (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[17102-:32] + (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[900-:32] - 1))) + 1)] = hpdcache_rsp_i[(hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1157-:32] * hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1285-:32]) + (hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32] + (hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1))-:(((hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1157-:32] * hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1285-:32]) + (hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32] + (hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1))) >= (hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32] + (hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 2)) ? (((hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1157-:32] * hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1285-:32]) + (hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32] + (hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1))) - (hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32] + (hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 2))) + 1 : ((hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32] + (hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 2)) - ((hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1157-:32] * hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1285-:32]) + (hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32] + (hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1)))) + 1)];
			// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:196:7
			assign cva6_req_o[dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[1124-:32] + (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[17102-:32] + (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[900-:32] - 1))-:((dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[1124-:32] + (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[17102-:32] + (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[900-:32] - 1))) >= (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[17102-:32] + (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[900-:32] + 0)) ? ((dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[1124-:32] + (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[17102-:32] + (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[900-:32] - 1))) - (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[17102-:32] + (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[900-:32] + 0))) + 1 : ((dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[17102-:32] + (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[900-:32] + 0)) - (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[1124-:32] + (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[17102-:32] + (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[900-:32] - 1)))) + 1)] = hpdcache_rsp_i[hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1-:((hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1) >= 2 ? hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 0 : 3 - (hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1))];
			// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:197:7
			assign cva6_req_o[2 + (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[1124-:32] + (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[17102-:32] + (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[900-:32] - 1)))] = hpdcache_req_ready_i;
			// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:199:7
			assign cva6_amo_resp_o[64] = hpdcache_rsp_valid_i && (hpdcache_rsp_i[hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1-:((hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1) >= 2 ? hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 0 : 3 - (hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1))] == {hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] {1'sb1}});
			// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:200:7
			assign cva6_amo_resp_o[63-:64] = (amo_is_word ? {{32 {amo_resp_word[31]}}, amo_resp_word} : hpdcache_rsp_i[((hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1157-:32] * hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1285-:32]) + (hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1093-:32] + (hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1125-:32] + 1))) - ((hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1157-:32] * hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1285-:32]) - 1)+:hpdcache_rsp_t_hpdcache_rsp_t_HPDcacheCfg[1285-:32]]);
			// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:204:7
			always @(posedge clk_i or negedge rst_ni) begin : amo_pending_ff
				// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:205:9
				if (!rst_ni)
					// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:206:11
					amo_pending_q <= 1'b0;
				else
					// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:208:11
					amo_pending_q <= ((cva6_amo_req_i[134] & hpdcache_req_ready_i) & ~amo_pending_q) | (~cva6_amo_resp_o[64] & amo_pending_q);
			end
		end
	endgenerate
	// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:221:3
	// removed an assertion item
	// forward_one_request_assert : assert property (@(posedge clk_i) 
	// 	$onehot0({forward_store, forward_amo})
	// ) else begin
	// 	// Trace: core/cache_subsystem/cva6_hpdcache_if_adapter.sv:223:8
	// 	$error("Only one request shall be forwarded");
	// end
	initial _sv2v_0 = 0;
endmodule
