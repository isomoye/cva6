module issue_read_operands_C2BA9_BE966 (
	clk_i,
	rst_ni,
	flush_i,
	stall_i,
	issue_instr_i,
	orig_instr_i,
	issue_instr_valid_i,
	issue_ack_o,
	rs1_o,
	rs1_i,
	rs1_valid_i,
	rs2_o,
	rs2_i,
	rs2_valid_i,
	rs3_o,
	rs3_i,
	rs3_valid_i,
	rd_clobber_gpr_i,
	rd_clobber_fpr_i,
	fu_data_o,
	rs1_forwarding_o,
	rs2_forwarding_o,
	pc_o,
	is_compressed_instr_o,
	flu_ready_i,
	alu_valid_o,
	branch_valid_o,
	tinst_o,
	branch_predict_o,
	lsu_ready_i,
	lsu_valid_o,
	mult_valid_o,
	fpu_ready_i,
	fpu_valid_o,
	fpu_fmt_o,
	fpu_rm_o,
	alu2_valid_o,
	csr_valid_o,
	cvxif_valid_o,
	cvxif_ready_i,
	cvxif_off_instr_o,
	hart_id_i,
	x_issue_ready_i,
	x_issue_resp_i,
	x_issue_valid_o,
	x_issue_req_o,
	x_register_ready_i,
	x_register_valid_o,
	x_register_o,
	x_commit_valid_o,
	x_commit_o,
	x_transaction_accepted_o,
	x_transaction_rejected_o,
	x_issue_writeback_o,
	x_id_o,
	waddr_i,
	wdata_i,
	we_gpr_i,
	we_fpr_i,
	stall_issue_o
);
	// removed localparam type branchpredict_sbe_t_branchpredict_sbe_t_CVA6Cfg_type
	parameter [17102:0] branchpredict_sbe_t_branchpredict_sbe_t_CVA6Cfg = 0;
	// removed localparam type fu_data_t_fu_data_t_CVA6Cfg_type
	parameter [17102:0] fu_data_t_fu_data_t_CVA6Cfg = 0;
	// removed localparam type rs3_len_t_CVA6Cfg_type
	parameter [17102:0] rs3_len_t_CVA6Cfg = 0;
	// removed localparam type scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg_type
	parameter [17102:0] scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg = 0;
	// removed localparam type x_commit_t_x_commit_t_x_commit_t_CVA6Cfg_type
	parameter [17102:0] x_commit_t_x_commit_t_x_commit_t_CVA6Cfg = 0;
	// removed localparam type x_issue_req_t_x_issue_req_t_x_issue_req_t_CVA6Cfg_type
	parameter [17102:0] x_issue_req_t_x_issue_req_t_x_issue_req_t_CVA6Cfg = 0;
	// removed localparam type x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg_type
	parameter [17102:0] x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg = 0;
	// removed localparam type x_register_t_x_register_t_x_register_t_CVA6Cfg_type
	parameter [17102:0] x_register_t_x_register_t_x_register_t_CVA6Cfg = 0;
	reg _sv2v_0;
	// removed import ariane_pkg::*;
	// Trace: core/issue_read_operands.sv:20:15
	localparam config_pkg_NrMaxRules = 16;
	// removed localparam type config_pkg_cache_type_t
	// removed localparam type config_pkg_noc_type_e
	// removed localparam type config_pkg_vm_mode_t
	// removed localparam type config_pkg_cva6_cfg_t
	localparam [17102:0] config_pkg_cva6_cfg_empty = 17103'd0;
	parameter [17102:0] CVA6Cfg = config_pkg_cva6_cfg_empty;
	// Trace: core/issue_read_operands.sv:21:20
	// removed localparam type branchpredict_sbe_t
	// Trace: core/issue_read_operands.sv:22:20
	// removed localparam type fu_data_t
	// Trace: core/issue_read_operands.sv:23:20
	// removed localparam type scoreboard_entry_t
	// Trace: core/issue_read_operands.sv:24:20
	// removed localparam type rs3_len_t
	// Trace: core/issue_read_operands.sv:25:20
	// removed localparam type x_issue_req_t
	// Trace: core/issue_read_operands.sv:26:20
	// removed localparam type x_issue_resp_t
	// Trace: core/issue_read_operands.sv:27:20
	// removed localparam type x_register_t
	// Trace: core/issue_read_operands.sv:28:20
	// removed localparam type x_commit_t
	// Trace: core/issue_read_operands.sv:32:5
	input wire clk_i;
	// Trace: core/issue_read_operands.sv:34:5
	input wire rst_ni;
	// Trace: core/issue_read_operands.sv:36:5
	input wire flush_i;
	// Trace: core/issue_read_operands.sv:38:5
	input wire stall_i;
	// Trace: core/issue_read_operands.sv:40:5
	input wire [((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (CVA6Cfg[16841-:32] * (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5)) - 1 : (CVA6Cfg[16841-:32] * (1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 3)):((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 0 : ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)] issue_instr_i;
	// Trace: core/issue_read_operands.sv:42:5
	input wire [(CVA6Cfg[16841-:32] * 32) - 1:0] orig_instr_i;
	// Trace: core/issue_read_operands.sv:44:5
	input wire [CVA6Cfg[16841-:32] - 1:0] issue_instr_valid_i;
	// Trace: core/issue_read_operands.sv:46:5
	output reg [CVA6Cfg[16841-:32] - 1:0] issue_ack_o;
	// Trace: core/issue_read_operands.sv:48:5
	localparam ariane_pkg_REG_ADDR_SIZE = 5;
	output reg [(CVA6Cfg[16841-:32] * 5) - 1:0] rs1_o;
	// Trace: core/issue_read_operands.sv:50:5
	input wire [(CVA6Cfg[16841-:32] * CVA6Cfg[17102-:32]) - 1:0] rs1_i;
	// Trace: core/issue_read_operands.sv:52:5
	input wire [CVA6Cfg[16841-:32] - 1:0] rs1_valid_i;
	// Trace: core/issue_read_operands.sv:54:5
	output reg [(CVA6Cfg[16841-:32] * 5) - 1:0] rs2_o;
	// Trace: core/issue_read_operands.sv:56:5
	input wire [(CVA6Cfg[16841-:32] * CVA6Cfg[17102-:32]) - 1:0] rs2_i;
	// Trace: core/issue_read_operands.sv:58:5
	input wire [CVA6Cfg[16841-:32] - 1:0] rs2_valid_i;
	// Trace: core/issue_read_operands.sv:60:5
	output reg [(CVA6Cfg[16841-:32] * 5) - 1:0] rs3_o;
	// Trace: core/issue_read_operands.sv:62:5
	input wire [(CVA6Cfg[16841-:32] * (rs3_len_t_CVA6Cfg[16433-:32] == 3 ? rs3_len_t_CVA6Cfg[17102-:32] : rs3_len_t_CVA6Cfg[16469-:32])) - 1:0] rs3_i;
	// Trace: core/issue_read_operands.sv:64:5
	input wire [CVA6Cfg[16841-:32] - 1:0] rs3_valid_i;
	// Trace: core/issue_read_operands.sv:67:5
	// removed localparam type ariane_pkg_fu_t
	input wire [127:0] rd_clobber_gpr_i;
	// Trace: core/issue_read_operands.sv:69:5
	input wire [127:0] rd_clobber_fpr_i;
	// Trace: core/issue_read_operands.sv:71:5
	output wire [(CVA6Cfg[16841-:32] * ((((12 + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[16503-:32])) - 1:0] fu_data_o;
	// Trace: core/issue_read_operands.sv:73:5
	output wire [(CVA6Cfg[16841-:32] * CVA6Cfg[17102-:32]) - 1:0] rs1_forwarding_o;
	// Trace: core/issue_read_operands.sv:75:5
	output wire [(CVA6Cfg[16841-:32] * CVA6Cfg[17102-:32]) - 1:0] rs2_forwarding_o;
	// Trace: core/issue_read_operands.sv:77:5
	output reg [CVA6Cfg[17070-:32] - 1:0] pc_o;
	// Trace: core/issue_read_operands.sv:79:5
	output reg is_compressed_instr_o;
	// Trace: core/issue_read_operands.sv:81:5
	input wire flu_ready_i;
	// Trace: core/issue_read_operands.sv:83:5
	output wire [CVA6Cfg[16841-:32] - 1:0] alu_valid_o;
	// Trace: core/issue_read_operands.sv:85:5
	output wire [CVA6Cfg[16841-:32] - 1:0] branch_valid_o;
	// Trace: core/issue_read_operands.sv:87:5
	output wire [(CVA6Cfg[16841-:32] * 32) - 1:0] tinst_o;
	// Trace: core/issue_read_operands.sv:89:5
	output reg [(3 + branchpredict_sbe_t_branchpredict_sbe_t_CVA6Cfg[17070-:32]) - 1:0] branch_predict_o;
	// Trace: core/issue_read_operands.sv:91:5
	input wire lsu_ready_i;
	// Trace: core/issue_read_operands.sv:93:5
	output wire [CVA6Cfg[16841-:32] - 1:0] lsu_valid_o;
	// Trace: core/issue_read_operands.sv:95:5
	output wire [CVA6Cfg[16841-:32] - 1:0] mult_valid_o;
	// Trace: core/issue_read_operands.sv:97:5
	input wire fpu_ready_i;
	// Trace: core/issue_read_operands.sv:99:5
	output wire [CVA6Cfg[16841-:32] - 1:0] fpu_valid_o;
	// Trace: core/issue_read_operands.sv:101:5
	output wire [1:0] fpu_fmt_o;
	// Trace: core/issue_read_operands.sv:103:5
	output wire [2:0] fpu_rm_o;
	// Trace: core/issue_read_operands.sv:105:5
	output wire [CVA6Cfg[16841-:32] - 1:0] alu2_valid_o;
	// Trace: core/issue_read_operands.sv:107:5
	output wire [CVA6Cfg[16841-:32] - 1:0] csr_valid_o;
	// Trace: core/issue_read_operands.sv:109:5
	output wire [CVA6Cfg[16841-:32] - 1:0] cvxif_valid_o;
	// Trace: core/issue_read_operands.sv:111:5
	input wire cvxif_ready_i;
	// Trace: core/issue_read_operands.sv:113:5
	output wire [31:0] cvxif_off_instr_o;
	// Trace: core/issue_read_operands.sv:115:5
	input wire [CVA6Cfg[17102-:32] - 1:0] hart_id_i;
	// Trace: core/issue_read_operands.sv:117:5
	input wire x_issue_ready_i;
	// Trace: core/issue_read_operands.sv:118:5
	input wire [((1 + (x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[63-:32] >= 0 ? x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[63-:32] + 1 : 1 - x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[63-:32])) + (x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[287-:32] + x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[95-:32])) - 1:0] x_issue_resp_i;
	// Trace: core/issue_read_operands.sv:119:5
	output wire x_issue_valid_o;
	// Trace: core/issue_read_operands.sv:120:5
	output wire [((32 + x_issue_req_t_x_issue_req_t_x_issue_req_t_CVA6Cfg[127-:32]) + x_issue_req_t_x_issue_req_t_x_issue_req_t_CVA6Cfg[255-:32]) - 1:0] x_issue_req_o;
	// Trace: core/issue_read_operands.sv:122:5
	input wire x_register_ready_i;
	// Trace: core/issue_read_operands.sv:123:5
	output wire x_register_valid_o;
	// Trace: core/issue_read_operands.sv:124:5
	output wire [(((x_register_t_x_register_t_x_register_t_CVA6Cfg[127-:32] + x_register_t_x_register_t_x_register_t_CVA6Cfg[255-:32]) + (x_register_t_x_register_t_x_register_t_CVA6Cfg[287-:32] * x_register_t_x_register_t_x_register_t_CVA6Cfg[223-:32])) + (x_register_t_x_register_t_x_register_t_CVA6Cfg[287-:32] + x_register_t_x_register_t_x_register_t_CVA6Cfg[95-:32])) - 1:0] x_register_o;
	// Trace: core/issue_read_operands.sv:126:5
	output wire x_commit_valid_o;
	// Trace: core/issue_read_operands.sv:127:5
	output wire [(x_commit_t_x_commit_t_x_commit_t_CVA6Cfg[127-:32] + x_commit_t_x_commit_t_x_commit_t_CVA6Cfg[255-:32]) + 0:0] x_commit_o;
	// Trace: core/issue_read_operands.sv:129:5
	output wire x_transaction_accepted_o;
	// Trace: core/issue_read_operands.sv:130:5
	output reg x_transaction_rejected_o;
	// Trace: core/issue_read_operands.sv:131:5
	output wire x_issue_writeback_o;
	// Trace: core/issue_read_operands.sv:132:5
	output wire [CVA6Cfg[16503-:32] - 1:0] x_id_o;
	// Trace: core/issue_read_operands.sv:134:5
	input wire [(CVA6Cfg[16873-:32] * 5) - 1:0] waddr_i;
	// Trace: core/issue_read_operands.sv:136:5
	input wire [(CVA6Cfg[16873-:32] * CVA6Cfg[17102-:32]) - 1:0] wdata_i;
	// Trace: core/issue_read_operands.sv:138:5
	input wire [CVA6Cfg[16873-:32] - 1:0] we_gpr_i;
	// Trace: core/issue_read_operands.sv:140:5
	input wire [CVA6Cfg[16873-:32] - 1:0] we_fpr_i;
	// Trace: core/issue_read_operands.sv:143:5
	output wire stall_issue_o;
	// Trace: core/issue_read_operands.sv:146:3
	localparam OPERANDS_PER_INSTR = CVA6Cfg[16433-:32] / CVA6Cfg[16841-:32];
	// Trace: core/issue_read_operands.sv:148:3
	// removed localparam type fus_busy_t
	// Trace: core/issue_read_operands.sv:152:3
	reg [CVA6Cfg[16841-:32] - 1:0] stall_raw;
	reg [CVA6Cfg[16841-:32] - 1:0] stall_waw;
	reg [CVA6Cfg[16841-:32] - 1:0] stall_rs1;
	reg [CVA6Cfg[16841-:32] - 1:0] stall_rs2;
	reg [CVA6Cfg[16841-:32] - 1:0] stall_rs3;
	// Trace: core/issue_read_operands.sv:153:3
	reg [CVA6Cfg[16841-:32] - 1:0] fu_busy;
	// Trace: core/issue_read_operands.sv:154:3
	reg [(CVA6Cfg[16841-:32] * 12) - 1:0] fus_busy;
	// Trace: core/issue_read_operands.sv:155:3
	reg [CVA6Cfg[16841-:32] - 1:0] issue_ack;
	// Trace: core/issue_read_operands.sv:157:3
	wire [(CVA6Cfg[16841-:32] * CVA6Cfg[17102-:32]) - 1:0] operand_a_regfile;
	wire [(CVA6Cfg[16841-:32] * CVA6Cfg[17102-:32]) - 1:0] operand_b_regfile;
	// Trace: core/issue_read_operands.sv:159:3
	wire [(CVA6Cfg[16841-:32] * (rs3_len_t_CVA6Cfg[16433-:32] == 3 ? rs3_len_t_CVA6Cfg[17102-:32] : rs3_len_t_CVA6Cfg[16469-:32])) - 1:0] operand_c_regfile;
	wire [(CVA6Cfg[16841-:32] * (rs3_len_t_CVA6Cfg[16433-:32] == 3 ? rs3_len_t_CVA6Cfg[17102-:32] : rs3_len_t_CVA6Cfg[16469-:32])) - 1:0] operand_c_gpr;
	// Trace: core/issue_read_operands.sv:160:3
	wire [(rs3_len_t_CVA6Cfg[16433-:32] == 3 ? rs3_len_t_CVA6Cfg[17102-:32] : rs3_len_t_CVA6Cfg[16469-:32]) - 1:0] operand_c_fpr;
	// Trace: core/issue_read_operands.sv:162:3
	reg [(CVA6Cfg[16841-:32] * ((((12 + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[16503-:32])) - 1:0] fu_data_n;
	reg [(CVA6Cfg[16841-:32] * ((((12 + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[16503-:32])) - 1:0] fu_data_q;
	// Trace: core/issue_read_operands.sv:163:3
	wire [CVA6Cfg[17102-:32] - 1:0] imm_forward_rs3;
	// Trace: core/issue_read_operands.sv:165:3
	reg [CVA6Cfg[16841-:32] - 1:0] alu_valid_q;
	// Trace: core/issue_read_operands.sv:166:3
	reg [CVA6Cfg[16841-:32] - 1:0] mult_valid_q;
	// Trace: core/issue_read_operands.sv:167:3
	reg [CVA6Cfg[16841-:32] - 1:0] fpu_valid_q;
	// Trace: core/issue_read_operands.sv:168:3
	reg [1:0] fpu_fmt_q;
	// Trace: core/issue_read_operands.sv:169:3
	reg [2:0] fpu_rm_q;
	// Trace: core/issue_read_operands.sv:170:3
	reg [CVA6Cfg[16841-:32] - 1:0] alu2_valid_q;
	// Trace: core/issue_read_operands.sv:171:3
	reg [CVA6Cfg[16841-:32] - 1:0] lsu_valid_q;
	// Trace: core/issue_read_operands.sv:172:3
	reg [CVA6Cfg[16841-:32] - 1:0] csr_valid_q;
	// Trace: core/issue_read_operands.sv:173:3
	reg [CVA6Cfg[16841-:32] - 1:0] branch_valid_q;
	// Trace: core/issue_read_operands.sv:174:3
	reg [CVA6Cfg[16841-:32] - 1:0] cvxif_valid_q;
	// Trace: core/issue_read_operands.sv:175:3
	reg [31:0] cvxif_off_instr_q;
	// Trace: core/issue_read_operands.sv:176:3
	wire cvxif_instruction_valid;
	// Trace: core/issue_read_operands.sv:179:3
	reg [(CVA6Cfg[16841-:32] * 32) - 1:0] tinst_n;
	reg [(CVA6Cfg[16841-:32] * 32) - 1:0] tinst_q;
	// Trace: core/issue_read_operands.sv:182:3
	reg [CVA6Cfg[16841-:32] - 1:0] forward_rs1;
	reg [CVA6Cfg[16841-:32] - 1:0] forward_rs2;
	reg [CVA6Cfg[16841-:32] - 1:0] forward_rs3;
	// Trace: core/issue_read_operands.sv:185:3
	// removed localparam type riscv_atype_t
	// removed localparam type riscv_itype_t
	// removed localparam type riscv_r4type_t
	// removed localparam type riscv_rftype_t
	// removed localparam type riscv_rtype_t
	// removed localparam type riscv_rvftype_t
	// removed localparam type riscv_stype_t
	// removed localparam type riscv_utype_t
	// removed localparam type riscv_instruction_t
	wire [31:0] orig_instr;
	// Trace: core/issue_read_operands.sv:186:3
	assign orig_instr = orig_instr_i[0+:32];
	// Trace: core/issue_read_operands.sv:189:3
	wire cvxif_req_allowed;
	// Trace: core/issue_read_operands.sv:190:3
	wire x_transaction_rejected;
	// Trace: core/issue_read_operands.sv:191:3
	wire [OPERANDS_PER_INSTR - 1:0] rs_valid;
	// Trace: core/issue_read_operands.sv:192:3
	wire [(OPERANDS_PER_INSTR * CVA6Cfg[17102-:32]) - 1:0] rs;
	// Trace: core/issue_read_operands.sv:194:3
	cvxif_issue_register_commit_if_driver_438A7_844C7 #(
		.x_commit_t_x_commit_t_x_commit_t_x_commit_t_CVA6Cfg(x_commit_t_x_commit_t_x_commit_t_CVA6Cfg),
		.x_issue_req_t_x_issue_req_t_x_issue_req_t_x_issue_req_t_CVA6Cfg(x_issue_req_t_x_issue_req_t_x_issue_req_t_CVA6Cfg),
		.x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg(x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg),
		.x_register_t_x_register_t_x_register_t_x_register_t_CVA6Cfg(x_register_t_x_register_t_x_register_t_CVA6Cfg),
		.CVA6Cfg(CVA6Cfg)
	) i_cvxif_issue_register_commit_if_driver(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(flush_i),
		.hart_id_i(hart_id_i),
		.issue_ready_i(x_issue_ready_i),
		.issue_resp_i(x_issue_resp_i),
		.issue_valid_o(x_issue_valid_o),
		.issue_req_o(x_issue_req_o),
		.register_ready_i(x_register_ready_i),
		.register_valid_o(x_register_valid_o),
		.register_o(x_register_o),
		.commit_valid_o(x_commit_valid_o),
		.commit_o(x_commit_o),
		.valid_i(cvxif_instruction_valid),
		.x_off_instr_i(orig_instr_i[0+:32]),
		.x_trans_id_i(issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 0 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) : ((0 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))))) + ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) >= (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + 1)) - 1)-:((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) >= (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + 1)]),
		.register_i(rs),
		.rs_valid_i(rs_valid),
		.cvxif_busy_o()
	);
	// Trace: core/issue_read_operands.sv:221:3
	generate
		if (OPERANDS_PER_INSTR == 3) begin : genblk1
			// Trace: core/issue_read_operands.sv:222:5
			assign rs_valid = {~stall_rs3[0], ~stall_rs2[0], ~stall_rs1[0]};
			// Trace: core/issue_read_operands.sv:223:5
			assign rs = {fu_data_n[0 + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1))-:((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1)) >= (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] + 0) ? ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1)) - (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] + 0)) + 1 : ((fu_data_t_fu_data_t_CVA6Cfg[16503-:32] + 0) - (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1))) + 1)], fu_data_n[0 + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1)))-:((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1))) >= (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] + 0)) ? ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1))) - (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] + 0))) + 1 : ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] + 0)) - (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1)))) + 1)], fu_data_n[0 + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1))))-:((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1)))) >= (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] + 0))) ? ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1)))) - (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] + 0)))) + 1 : ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] + 0))) - (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1))))) + 1)]};
		end
		else begin : genblk1
			// Trace: core/issue_read_operands.sv:225:5
			assign rs_valid = {~stall_rs2[0], ~stall_rs1[0]};
			// Trace: core/issue_read_operands.sv:226:5
			assign rs = {fu_data_n[0 + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1)))-:((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1))) >= (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] + 0)) ? ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1))) - (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] + 0))) + 1 : ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] + 0)) - (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1)))) + 1)], fu_data_n[0 + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1))))-:((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1)))) >= (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] + 0))) ? ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1)))) - (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] + 0)))) + 1 : ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] + 0))) - (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1))))) + 1)]};
		end
	endgenerate
	// Trace: core/issue_read_operands.sv:231:3
	assign cvxif_req_allowed = (issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 0 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : ((0 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] == 4'd9) && !stall_waw[0];
	// Trace: core/issue_read_operands.sv:232:3
	assign cvxif_instruction_valid = (!issue_instr_i[0 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) : (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) : (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))] && issue_instr_valid_i[0]) && cvxif_req_allowed;
	// Trace: core/issue_read_operands.sv:233:3
	assign x_transaction_accepted_o = (x_issue_valid_o && x_issue_ready_i) && x_issue_resp_i[1 + ((x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[63-:32] >= 0 ? x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[63-:32] + 1 : 1 - x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[63-:32]) + ((x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[287-:32] + x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[95-:32]) - 1))];
	// Trace: core/issue_read_operands.sv:234:3
	assign x_transaction_rejected = (x_issue_valid_o && x_issue_ready_i) && ~x_issue_resp_i[1 + ((x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[63-:32] >= 0 ? x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[63-:32] + 1 : 1 - x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[63-:32]) + ((x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[287-:32] + x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[95-:32]) - 1))];
	// Trace: core/issue_read_operands.sv:235:3
	assign x_issue_writeback_o = x_issue_resp_i[(x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[63-:32] >= 0 ? x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[63-:32] + 1 : 1 - x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[63-:32]) + ((x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[287-:32] + x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[95-:32]) - 1)-:(((x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[63-:32] >= 0 ? x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[63-:32] + 1 : 1 - x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[63-:32]) + ((x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[287-:32] + x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[95-:32]) - 1)) >= ((x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[287-:32] + x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[95-:32]) + 0) ? (((x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[63-:32] >= 0 ? x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[63-:32] + 1 : 1 - x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[63-:32]) + ((x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[287-:32] + x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[95-:32]) - 1)) - ((x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[287-:32] + x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[95-:32]) + 0)) + 1 : (((x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[287-:32] + x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[95-:32]) + 0) - ((x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[63-:32] >= 0 ? x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[63-:32] + 1 : 1 - x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[63-:32]) + ((x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[287-:32] + x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[95-:32]) - 1))) + 1)];
	// Trace: core/issue_read_operands.sv:236:3
	assign x_id_o = x_issue_req_o[x_issue_req_t_x_issue_req_t_x_issue_req_t_CVA6Cfg[255-:32] - 1-:x_issue_req_t_x_issue_req_t_x_issue_req_t_CVA6Cfg[255-:32]];
	// Trace: core/issue_read_operands.sv:240:3
	genvar _gv_i_34;
	generate
		for (_gv_i_34 = 0; _gv_i_34 < CVA6Cfg[16841-:32]; _gv_i_34 = _gv_i_34 + 1) begin : genblk2
			localparam i = _gv_i_34;
			// Trace: core/issue_read_operands.sv:241:5
			assign rs1_forwarding_o[i * CVA6Cfg[17102-:32]+:CVA6Cfg[17102-:32]] = fu_data_n[(i * ((((12 + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[16503-:32])) + (((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1)))) - ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] - 1) - (CVA6Cfg[17070-:32] - 1))) >= ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1)))) - (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] - 1)) ? (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1)))) - ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] - 1) - (CVA6Cfg[17070-:32] - 1)) : (((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1)))) - ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] - 1) - (CVA6Cfg[17070-:32] - 1))) + (((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1)))) - ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] - 1) - (CVA6Cfg[17070-:32] - 1))) >= ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1)))) - (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] - 1)) ? (((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1)))) - ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] - 1) - (CVA6Cfg[17070-:32] - 1))) - ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1)))) - (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] - 1))) + 1 : (((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1)))) - (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] - 1)) - ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1)))) - ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] - 1) - (CVA6Cfg[17070-:32] - 1)))) + 1)) - 1)-:(((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1)))) - ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] - 1) - (CVA6Cfg[17070-:32] - 1))) >= ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1)))) - (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] - 1)) ? (((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1)))) - ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] - 1) - (CVA6Cfg[17070-:32] - 1))) - ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1)))) - (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] - 1))) + 1 : (((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1)))) - (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] - 1)) - ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1)))) - ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] - 1) - (CVA6Cfg[17070-:32] - 1)))) + 1)];
			// Trace: core/issue_read_operands.sv:242:5
			assign rs2_forwarding_o[i * CVA6Cfg[17102-:32]+:CVA6Cfg[17102-:32]] = fu_data_n[(i * ((((12 + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[16503-:32])) + (((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1))) - ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] - 1) - (CVA6Cfg[17070-:32] - 1))) >= ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1))) - (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] - 1)) ? (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1))) - ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] - 1) - (CVA6Cfg[17070-:32] - 1)) : (((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1))) - ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] - 1) - (CVA6Cfg[17070-:32] - 1))) + (((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1))) - ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] - 1) - (CVA6Cfg[17070-:32] - 1))) >= ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1))) - (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] - 1)) ? (((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1))) - ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] - 1) - (CVA6Cfg[17070-:32] - 1))) - ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1))) - (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] - 1))) + 1 : (((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1))) - (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] - 1)) - ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1))) - ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] - 1) - (CVA6Cfg[17070-:32] - 1)))) + 1)) - 1)-:(((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1))) - ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] - 1) - (CVA6Cfg[17070-:32] - 1))) >= ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1))) - (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] - 1)) ? (((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1))) - ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] - 1) - (CVA6Cfg[17070-:32] - 1))) - ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1))) - (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] - 1))) + 1 : (((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1))) - (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] - 1)) - ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1))) - ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] - 1) - (CVA6Cfg[17070-:32] - 1)))) + 1)];
		end
	endgenerate
	// Trace: core/issue_read_operands.sv:245:3
	assign fu_data_o = fu_data_q;
	// Trace: core/issue_read_operands.sv:246:3
	assign alu_valid_o = alu_valid_q;
	// Trace: core/issue_read_operands.sv:247:3
	assign branch_valid_o = branch_valid_q;
	// Trace: core/issue_read_operands.sv:248:3
	assign lsu_valid_o = lsu_valid_q;
	// Trace: core/issue_read_operands.sv:249:3
	assign csr_valid_o = csr_valid_q;
	// Trace: core/issue_read_operands.sv:250:3
	assign mult_valid_o = mult_valid_q;
	// Trace: core/issue_read_operands.sv:251:3
	assign fpu_valid_o = fpu_valid_q;
	// Trace: core/issue_read_operands.sv:252:3
	assign fpu_fmt_o = fpu_fmt_q;
	// Trace: core/issue_read_operands.sv:253:3
	assign fpu_rm_o = fpu_rm_q;
	// Trace: core/issue_read_operands.sv:254:3
	assign alu2_valid_o = alu2_valid_q;
	// Trace: core/issue_read_operands.sv:255:3
	assign cvxif_valid_o = (CVA6Cfg[16539] ? cvxif_valid_q : {CVA6Cfg[16841-:32] {1'sb0}});
	// Trace: core/issue_read_operands.sv:256:3
	assign cvxif_off_instr_o = (CVA6Cfg[16539] ? cvxif_off_instr_q : {32 {1'sb0}});
	// Trace: core/issue_read_operands.sv:257:3
	assign stall_issue_o = stall_raw[0];
	// Trace: core/issue_read_operands.sv:258:3
	assign tinst_o = (CVA6Cfg[16543] ? tinst_q : {CVA6Cfg[16841-:32] * 32 {1'sb0}});
	// Trace: core/issue_read_operands.sv:263:3
	// removed localparam type ariane_pkg_fu_op
	always @(*) begin : structural_hazards
		if (_sv2v_0)
			;
		// Trace: core/issue_read_operands.sv:264:5
		fus_busy = 1'sb0;
		// Trace: core/issue_read_operands.sv:268:5
		if (!flu_ready_i) begin
			// Trace: core/issue_read_operands.sv:269:7
			fus_busy[8] = 1'b1;
			// Trace: core/issue_read_operands.sv:270:7
			fus_busy[6] = 1'b1;
			// Trace: core/issue_read_operands.sv:271:7
			fus_busy[4] = 1'b1;
			// Trace: core/issue_read_operands.sv:272:7
			fus_busy[5] = 1'b1;
		end
		if (mult_valid_q) begin
			// Trace: core/issue_read_operands.sv:278:7
			fus_busy[8] = 1'b1;
			// Trace: core/issue_read_operands.sv:279:7
			fus_busy[6] = 1'b1;
			// Trace: core/issue_read_operands.sv:280:7
			fus_busy[4] = 1'b1;
		end
		if (CVA6Cfg[16471] && !fpu_ready_i) begin
			// Trace: core/issue_read_operands.sv:284:7
			fus_busy[3] = 1'b1;
			// Trace: core/issue_read_operands.sv:285:7
			fus_busy[2] = 1'b1;
			// Trace: core/issue_read_operands.sv:286:7
			if (CVA6Cfg[16874])
				// Trace: core/issue_read_operands.sv:286:34
				fus_busy[7] = 1'b1;
		end
		if (!lsu_ready_i) begin
			// Trace: core/issue_read_operands.sv:290:7
			fus_busy[10] = 1'b1;
			// Trace: core/issue_read_operands.sv:291:7
			fus_busy[9] = 1'b1;
		end
		if (CVA6Cfg[16874]) begin
			// Trace: core/issue_read_operands.sv:295:7
			fus_busy[12+:12] = fus_busy[0+:12];
			// Trace: core/issue_read_operands.sv:298:7
			fus_busy[16] = 1'b1;
			// Trace: core/issue_read_operands.sv:300:7
			fus_busy[13] = 1'b1;
			// Trace: core/issue_read_operands.sv:302:7
			(* full_case, parallel_case *)
			case (issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 0 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : ((0 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)])
				4'd0:
					// Trace: core/issue_read_operands.sv:303:16
					fus_busy[23] = 1'b1;
				4'd4:
					// Trace: core/issue_read_operands.sv:305:11
					if (CVA6Cfg[16809]) begin
						// Trace: core/issue_read_operands.sv:307:13
						fus_busy[20] = 1'b1;
						// Trace: core/issue_read_operands.sv:308:13
						fus_busy[18] = 1'b1;
						// Trace: core/issue_read_operands.sv:309:13
						fus_busy[16] = 1'b1;
						// Trace: core/issue_read_operands.sv:311:13
						fus_busy[22] = 1'b1;
						// Trace: core/issue_read_operands.sv:313:13
						fus_busy[21] = 1'b1;
					end
					else
						// Trace: core/issue_read_operands.sv:316:13
						if (issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 0 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : ((0 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] == 8'd0) begin
							// Trace: core/issue_read_operands.sv:317:15
							fus_busy[20] = 1'b1;
							// Trace: core/issue_read_operands.sv:318:15
							fus_busy[18] = 1'b1;
							// Trace: core/issue_read_operands.sv:319:15
							fus_busy[16] = 1'b1;
						end
						else
							// Trace: core/issue_read_operands.sv:322:15
							fus_busy[12+:12] = 1'sb1;
				4'd3:
					// Trace: core/issue_read_operands.sv:327:11
					if (CVA6Cfg[16874] && !fus_busy[7]) begin
						// Trace: core/issue_read_operands.sv:328:13
						fus_busy[19] = 1'b1;
						// Trace: core/issue_read_operands.sv:331:13
						fus_busy[15] = 1'b1;
						// Trace: core/issue_read_operands.sv:332:13
						fus_busy[14] = 1'b1;
					end
					else begin
						// Trace: core/issue_read_operands.sv:334:13
						fus_busy[20] = 1'b1;
						// Trace: core/issue_read_operands.sv:335:13
						fus_busy[18] = 1'b1;
						// Trace: core/issue_read_operands.sv:336:13
						fus_busy[16] = 1'b1;
					end
				4'd6:
					// Trace: core/issue_read_operands.sv:341:11
					fus_busy[12+:12] = 1'sb1;
				4'd5:
					// Trace: core/issue_read_operands.sv:343:16
					fus_busy[17] = 1'b1;
				4'd7, 4'd8: begin
					// Trace: core/issue_read_operands.sv:345:11
					fus_busy[15] = 1'b1;
					// Trace: core/issue_read_operands.sv:346:11
					fus_busy[14] = 1'b1;
				end
				4'd1, 4'd2: begin
					// Trace: core/issue_read_operands.sv:349:11
					fus_busy[22] = 1'b1;
					// Trace: core/issue_read_operands.sv:350:11
					fus_busy[21] = 1'b1;
				end
				4'd9:
					;
			endcase
		end
	end
	// Trace: core/issue_read_operands.sv:359:3
	genvar _gv_i_35;
	generate
		for (_gv_i_35 = 0; _gv_i_35 < CVA6Cfg[16841-:32]; _gv_i_35 = _gv_i_35 + 1) begin : genblk3
			localparam i = _gv_i_35;
			// Trace: core/issue_read_operands.sv:360:5
			always @(*) begin
				if (_sv2v_0)
					;
				// Trace: core/issue_read_operands.sv:361:7
				(* full_case, parallel_case *)
				case (issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)])
					4'd0:
						// Trace: core/issue_read_operands.sv:362:15
						fu_busy[i] = fus_busy[(i * 12) + 11];
					4'd3:
						// Trace: core/issue_read_operands.sv:364:11
						if (CVA6Cfg[16874] && !fus_busy[(i * 12) + 7])
							// Trace: core/issue_read_operands.sv:365:13
							fu_busy[i] = fus_busy[(i * 12) + 7];
						else
							// Trace: core/issue_read_operands.sv:367:13
							fu_busy[i] = fus_busy[(i * 12) + 8];
					4'd4:
						// Trace: core/issue_read_operands.sv:370:20
						fu_busy[i] = fus_busy[(i * 12) + 6];
					4'd6:
						// Trace: core/issue_read_operands.sv:371:14
						fu_busy[i] = fus_busy[(i * 12) + 4];
					4'd5:
						// Trace: core/issue_read_operands.sv:372:15
						fu_busy[i] = fus_busy[(i * 12) + 5];
					4'd1:
						// Trace: core/issue_read_operands.sv:373:15
						fu_busy[i] = fus_busy[(i * 12) + 10];
					4'd2:
						// Trace: core/issue_read_operands.sv:374:16
						fu_busy[i] = fus_busy[(i * 12) + 9];
					4'd9:
						// Trace: core/issue_read_operands.sv:375:16
						fu_busy[i] = fus_busy[(i * 12) + 1];
					default:
						if (CVA6Cfg[16471])
							// Trace: core/issue_read_operands.sv:378:11
							(* full_case, parallel_case *)
							case (issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)])
								4'd7:
									// Trace: core/issue_read_operands.sv:379:18
									fu_busy[i] = fus_busy[(i * 12) + 3];
								4'd8:
									// Trace: core/issue_read_operands.sv:380:22
									fu_busy[i] = fus_busy[(i * 12) + 2];
								default:
									// Trace: core/issue_read_operands.sv:381:22
									fu_busy[i] = 1'b0;
							endcase
						else
							// Trace: core/issue_read_operands.sv:384:11
							fu_busy[i] = 1'b0;
				endcase
			end
		end
	endgenerate
	// Trace: core/issue_read_operands.sv:395:3
	function automatic ariane_pkg_is_imm_fpr;
		// Trace: core/include/ariane_pkg.sv:578:39
		input reg [7:0] op;
		// Trace: core/include/ariane_pkg.sv:579:5
		(* full_case, parallel_case *)
		case (op)
			8'd104, 8'd105, 8'd110, 8'd111, 8'd112, 8'd113, 8'd133, 8'd134, 8'd135, 8'd136: ariane_pkg_is_imm_fpr = 1'b1;
			default: ariane_pkg_is_imm_fpr = 1'b0;
		endcase
	endfunction
	function automatic ariane_pkg_is_rd_fpr;
		// Trace: core/include/ariane_pkg.sv:597:38
		input reg [7:0] op;
		// Trace: core/include/ariane_pkg.sv:598:5
		(* full_case, parallel_case *)
		case (op)
			8'd96, 8'd97, 8'd98, 8'd99, 8'd104, 8'd105, 8'd106, 8'd107, 8'd108, 8'd109, 8'd110, 8'd111, 8'd112, 8'd113, 8'd115, 8'd116, 8'd117, 8'd119, 8'd122, 8'd123, 8'd124, 8'd125, 8'd126, 8'd133, 8'd134, 8'd135, 8'd136, 8'd183: ariane_pkg_is_rd_fpr = 1'b1;
			default: ariane_pkg_is_rd_fpr = 1'b0;
		endcase
	endfunction
	function automatic ariane_pkg_is_rs1_fpr;
		// Trace: core/include/ariane_pkg.sv:507:39
		input reg [7:0] op;
		// Trace: core/include/ariane_pkg.sv:508:5
		(* full_case, parallel_case *)
		case (op)
			8'd106, 8'd107, 8'd108, 8'd109, 8'd110, 8'd111, 8'd112, 8'd113, 8'd114, 8'd116, 8'd117, 8'd118, 8'd120, 8'd121, 8'd122, 8'd123, 8'd124, 8'd125, 8'd126, 8'd127, 8'd128, 8'd129, 8'd130, 8'd131, 8'd132, 8'd133, 8'd134, 8'd135, 8'd136, 8'd182: ariane_pkg_is_rs1_fpr = 1'b1;
			default: ariane_pkg_is_rs1_fpr = 1'b0;
		endcase
	endfunction
	function automatic ariane_pkg_is_rs2_fpr;
		// Trace: core/include/ariane_pkg.sv:546:39
		input reg [7:0] op;
		// Trace: core/include/ariane_pkg.sv:547:5
		(* full_case, parallel_case *)
		case (op)
			8'd100, 8'd101, 8'd102, 8'd103, 8'd104, 8'd105, 8'd106, 8'd107, 8'd108, 8'd110, 8'd111, 8'd112, 8'd113, 8'd116, 8'd117, 8'd118, 8'd120, 8'd122, 8'd123, 8'd124, 8'd125, 8'd126: ariane_pkg_is_rs2_fpr = 1'b1;
			default: ariane_pkg_is_rs2_fpr = 1'b0;
		endcase
	endfunction
	always @(*) begin : operands_available
		if (_sv2v_0)
			;
		// Trace: core/issue_read_operands.sv:396:5
		stall_raw = {CVA6Cfg[16841-:32] {stall_i}};
		// Trace: core/issue_read_operands.sv:397:5
		stall_rs1 = {CVA6Cfg[16841-:32] {stall_i}};
		// Trace: core/issue_read_operands.sv:398:5
		stall_rs2 = {CVA6Cfg[16841-:32] {stall_i}};
		// Trace: core/issue_read_operands.sv:399:5
		stall_rs3 = {CVA6Cfg[16841-:32] {stall_i}};
		// Trace: core/issue_read_operands.sv:401:5
		forward_rs1 = 1'sb0;
		// Trace: core/issue_read_operands.sv:402:5
		forward_rs2 = 1'sb0;
		// Trace: core/issue_read_operands.sv:403:5
		forward_rs3 = 1'sb0;
		// Trace: core/issue_read_operands.sv:405:5
		begin : sv2v_autoblock_1
			// Trace: core/issue_read_operands.sv:405:10
			reg [31:0] i;
			// Trace: core/issue_read_operands.sv:405:10
			for (i = 0; i < CVA6Cfg[16841-:32]; i = i + 1)
				begin
					// Trace: core/issue_read_operands.sv:407:7
					rs1_o[i * 5+:5] = issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)];
					// Trace: core/issue_read_operands.sv:408:7
					rs2_o[i * 5+:5] = issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)];
					// Trace: core/issue_read_operands.sv:409:7
					rs3_o[i * 5+:5] = issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5) : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) + (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1))) + 1 : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5))) + 1)) - 1) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5) : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) + (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1))) + 1 : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5))) + 1)) - 1)) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5) : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) + (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1))) + 1 : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5))) + 1)) - 1) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5) : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) + (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1))) + 1 : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5))) + 1)) - 1))) + (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1))) + 1 : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5))) + 1)) - 1)-:(((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1))) + 1 : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5))) + 1)];
					// Trace: core/issue_read_operands.sv:416:7
					if (!issue_instr_i[(i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 2 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (2 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))] && (CVA6Cfg[16471] && ariane_pkg_is_rs1_fpr(issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)]) ? rd_clobber_fpr_i[issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] * 4+:4] != 4'd0 : rd_clobber_gpr_i[issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] * 4+:4] != 4'd0)) begin
						begin
							// Trace: core/issue_read_operands.sv:423:9
							if (rs1_valid_i[i] && (CVA6Cfg[16471] && ariane_pkg_is_rs1_fpr(issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)]) ? 1'b1 : (rd_clobber_gpr_i[issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] * 4+:4] != 4'd6) || (CVA6Cfg[16366] && (issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] == 8'd30))))
								// Trace: core/issue_read_operands.sv:427:11
								forward_rs1[i] = 1'b1;
							else begin
								// Trace: core/issue_read_operands.sv:429:11
								stall_raw[i] = 1'b1;
								// Trace: core/issue_read_operands.sv:430:11
								stall_rs1[i] = 1'b1;
							end
						end
					end
					if ((CVA6Cfg[16471] && ariane_pkg_is_rs2_fpr(issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)]) ? rd_clobber_fpr_i[issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] * 4+:4] != 4'd0 : rd_clobber_gpr_i[issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] * 4+:4] != 4'd0)) begin
						begin
							// Trace: core/issue_read_operands.sv:439:9
							if (rs2_valid_i[i] && (CVA6Cfg[16471] && ariane_pkg_is_rs2_fpr(issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)]) ? 1'b1 : (rd_clobber_gpr_i[issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] * 4+:4] != 4'd6) || (CVA6Cfg[16366] && (issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] == 8'd30))))
								// Trace: core/issue_read_operands.sv:443:11
								forward_rs2[i] = 1'b1;
							else begin
								// Trace: core/issue_read_operands.sv:445:11
								stall_raw[i] = 1'b1;
								// Trace: core/issue_read_operands.sv:446:11
								stall_rs2[i] = 1'b1;
							end
						end
					end
					if ((CVA6Cfg[16471] && ariane_pkg_is_imm_fpr(issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)]) ? rd_clobber_fpr_i[issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5) : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) + (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1))) + 1 : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5))) + 1)) - 1) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5) : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) + (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1))) + 1 : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5))) + 1)) - 1)) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5) : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) + (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1))) + 1 : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5))) + 1)) - 1) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5) : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) + (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1))) + 1 : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5))) + 1)) - 1))) + (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1))) + 1 : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5))) + 1)) - 1)-:(((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1))) + 1 : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5))) + 1)] * 4+:4] != 4'd0 : 0)) begin
						begin
							// Trace: core/issue_read_operands.sv:455:9
							if (rs3_valid_i[i])
								// Trace: core/issue_read_operands.sv:456:11
								forward_rs3[i] = 1'b1;
							else begin
								// Trace: core/issue_read_operands.sv:458:11
								stall_raw[i] = 1'b1;
								// Trace: core/issue_read_operands.sv:459:11
								stall_rs3[i] = 1'b1;
							end
						end
					end
				end
		end
		if (CVA6Cfg[16539]) begin
			// Trace: core/issue_read_operands.sv:465:7
			if (x_issue_valid_o && x_issue_resp_i[1 + ((x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[63-:32] >= 0 ? x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[63-:32] + 1 : 1 - x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[63-:32]) + ((x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[287-:32] + x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[95-:32]) - 1))]) begin
				// Trace: core/issue_read_operands.sv:466:9
				if (~x_issue_resp_i[((x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[287-:32] + x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[95-:32]) - 1) - ((x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[287-:32] + x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[95-:32]) - 1)]) begin
					// Trace: core/issue_read_operands.sv:467:11
					forward_rs1[0] = 1'b0;
					// Trace: core/issue_read_operands.sv:468:11
					stall_rs1[0] = 1'b0;
				end
				if (~x_issue_resp_i[((x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[287-:32] + x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[95-:32]) - 1) - ((x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[287-:32] + x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[95-:32]) - 2)]) begin
					// Trace: core/issue_read_operands.sv:471:11
					forward_rs2[0] = 1'b0;
					// Trace: core/issue_read_operands.sv:472:11
					stall_rs2[0] = 1'b0;
				end
				if ((OPERANDS_PER_INSTR == 3) && ~x_issue_resp_i[((x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[287-:32] + x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[95-:32]) - 1) - ((x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[287-:32] + x_issue_resp_t_x_issue_resp_t_x_issue_resp_t_CVA6Cfg[95-:32]) - 3)]) begin
					// Trace: core/issue_read_operands.sv:475:11
					forward_rs3[0] = 1'b0;
					// Trace: core/issue_read_operands.sv:476:11
					stall_rs3[0] = 1'b0;
				end
			end
			// Trace: core/issue_read_operands.sv:479:7
			stall_raw[0] = (stall_rs1[0] || stall_rs2[0]) || stall_rs3[0];
		end
		if (CVA6Cfg[16874]) begin
			// Trace: core/issue_read_operands.sv:483:7
			if (((!issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 2 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (2 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))] && (!CVA6Cfg[16471] || (ariane_pkg_is_rs1_fpr(issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : ((((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)]) == ariane_pkg_is_rd_fpr(issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 0 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : ((0 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)])))) && (issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : ((((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] == issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 0 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : ((0 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)])) && (issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : ((((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] != {5 {1'sb0}}))
				// Trace: core/issue_read_operands.sv:488:9
				stall_raw[1] = 1'b1;
			if (((!CVA6Cfg[16471] || (ariane_pkg_is_rs2_fpr(issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : ((((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)]) == ariane_pkg_is_rd_fpr(issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 0 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : ((0 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)]))) && (issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : ((((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] == issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 0 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : ((0 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)])) && (issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : ((((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] != {5 {1'sb0}}))
				// Trace: core/issue_read_operands.sv:496:9
				stall_raw[1] = 1'b1;
			if ((CVA6Cfg[16471] && ariane_pkg_is_imm_fpr(issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : ((((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)]) ? ariane_pkg_is_rd_fpr(issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 0 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : ((0 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)]) && (issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 0 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : ((0 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] == issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5) : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) + (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1))) + 1 : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5))) + 1)) - 1) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5) : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) + (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1))) + 1 : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5))) + 1)) - 1)) : ((((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5) : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) + (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1))) + 1 : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5))) + 1)) - 1) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5) : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) + (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1))) + 1 : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5))) + 1)) - 1))) + (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1))) + 1 : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5))) + 1)) - 1)-:(((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1))) + 1 : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5))) + 1)]) : ((issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : ((((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] == 8'd137) && (OPERANDS_PER_INSTR == 3) ? issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 0 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : ((0 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] == issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5) : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) + (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1))) + 1 : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5))) + 1)) - 1) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5) : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) + (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1))) + 1 : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5))) + 1)) - 1)) : ((((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5) : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) + (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1))) + 1 : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5))) + 1)) - 1) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5) : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) + (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1))) + 1 : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5))) + 1)) - 1))) + (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1))) + 1 : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5))) + 1)) - 1)-:(((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1))) + 1 : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5))) + 1)] : 1'b0)))
				// Trace: core/issue_read_operands.sv:507:9
				stall_raw[1] = 1'b1;
		end
	end
	// Trace: core/issue_read_operands.sv:513:3
	generate
		if (OPERANDS_PER_INSTR == 3) begin : gen_gp_rs3
			// Trace: core/issue_read_operands.sv:514:5
			assign imm_forward_rs3 = rs3_i[0+:(rs3_len_t_CVA6Cfg[16433-:32] == 3 ? rs3_len_t_CVA6Cfg[17102-:32] : rs3_len_t_CVA6Cfg[16469-:32])];
		end
		else begin : gen_fp_rs3
			// Trace: core/issue_read_operands.sv:516:5
			assign imm_forward_rs3 = {{CVA6Cfg[17102-:32] - CVA6Cfg[16469-:32] {1'b0}}, rs3_i[0+:(rs3_len_t_CVA6Cfg[16433-:32] == 3 ? rs3_len_t_CVA6Cfg[17102-:32] : rs3_len_t_CVA6Cfg[16469-:32])]};
		end
	endgenerate
	// Trace: core/issue_read_operands.sv:520:3
	genvar _gv_i_36;
	generate
		for (_gv_i_36 = 0; _gv_i_36 < CVA6Cfg[16841-:32]; _gv_i_36 = _gv_i_36 + 1) begin : genblk5
			localparam i = _gv_i_36;
			// Trace: core/issue_read_operands.sv:521:5
			always @(*) begin : forwarding_operand_select
				if (_sv2v_0)
					;
				// Trace: core/issue_read_operands.sv:523:7
				fu_data_n[(i * ((((12 + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[16503-:32])) + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1))))-:((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1)))) >= (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] + 0))) ? ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1)))) - (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] + 0)))) + 1 : ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] + 0))) - (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1))))) + 1)] = operand_a_regfile[i * CVA6Cfg[17102-:32]+:CVA6Cfg[17102-:32]];
				// Trace: core/issue_read_operands.sv:524:7
				fu_data_n[(i * ((((12 + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[16503-:32])) + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1)))-:((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1))) >= (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] + 0)) ? ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1))) - (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] + 0))) + 1 : ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] + 0)) - (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1)))) + 1)] = operand_b_regfile[i * CVA6Cfg[17102-:32]+:CVA6Cfg[17102-:32]];
				// Trace: core/issue_read_operands.sv:528:7
				if (OPERANDS_PER_INSTR == 3)
					// Trace: core/issue_read_operands.sv:529:9
					fu_data_n[(i * ((((12 + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[16503-:32])) + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1))-:((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1)) >= (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] + 0) ? ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1)) - (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] + 0)) + 1 : ((fu_data_t_fu_data_t_CVA6Cfg[16503-:32] + 0) - (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1))) + 1)] = (CVA6Cfg[16471] && ariane_pkg_is_imm_fpr(issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)]) ? {{CVA6Cfg[17102-:32] - CVA6Cfg[16469-:32] {1'b0}}, operand_c_regfile[i * (rs3_len_t_CVA6Cfg[16433-:32] == 3 ? rs3_len_t_CVA6Cfg[17102-:32] : rs3_len_t_CVA6Cfg[16469-:32])+:(rs3_len_t_CVA6Cfg[16433-:32] == 3 ? rs3_len_t_CVA6Cfg[17102-:32] : rs3_len_t_CVA6Cfg[16469-:32])]} : (issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] == 8'd137 ? operand_c_regfile[i * (rs3_len_t_CVA6Cfg[16433-:32] == 3 ? rs3_len_t_CVA6Cfg[17102-:32] : rs3_len_t_CVA6Cfg[16469-:32])+:(rs3_len_t_CVA6Cfg[16433-:32] == 3 ? rs3_len_t_CVA6Cfg[17102-:32] : rs3_len_t_CVA6Cfg[16469-:32])] : issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) >= (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) + 1 : ((4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + 1)) - 1)-:((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) >= (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) + 1 : ((4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + 1)]));
				else
					// Trace: core/issue_read_operands.sv:533:9
					fu_data_n[(i * ((((12 + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[16503-:32])) + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1))-:((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1)) >= (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] + 0) ? ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1)) - (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] + 0)) + 1 : ((fu_data_t_fu_data_t_CVA6Cfg[16503-:32] + 0) - (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1))) + 1)] = (CVA6Cfg[16471] && ariane_pkg_is_imm_fpr(issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)]) ? {{CVA6Cfg[17102-:32] - CVA6Cfg[16469-:32] {1'b0}}, operand_c_regfile[i * (rs3_len_t_CVA6Cfg[16433-:32] == 3 ? rs3_len_t_CVA6Cfg[17102-:32] : rs3_len_t_CVA6Cfg[16469-:32])+:(rs3_len_t_CVA6Cfg[16433-:32] == 3 ? rs3_len_t_CVA6Cfg[17102-:32] : rs3_len_t_CVA6Cfg[16469-:32])]} : issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) >= (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) + 1 : ((4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + 1)) - 1)-:((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) >= (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) + 1 : ((4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + 1)]);
				// Trace: core/issue_read_operands.sv:536:7
				fu_data_n[(i * ((((12 + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[16503-:32])) + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1)-:fu_data_t_fu_data_t_CVA6Cfg[16503-:32]] = issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))))) + ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) >= (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + 1)) - 1)-:((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) >= (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + 1)];
				// Trace: core/issue_read_operands.sv:537:7
				fu_data_n[(i * ((((12 + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[16503-:32])) + (12 + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1)))))-:((12 + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1))))) >= (8 + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] + 0))))) ? ((12 + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1))))) - (8 + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] + 0)))))) + 1 : ((8 + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] + 0))))) - (12 + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1)))))) + 1)] = issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)];
				// Trace: core/issue_read_operands.sv:538:7
				fu_data_n[(i * ((((12 + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[16503-:32])) + (8 + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1)))))-:((8 + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1))))) >= (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] + 0)))) ? ((8 + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1))))) - (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] + 0))))) + 1 : ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] + 0)))) - (8 + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1)))))) + 1)] = issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)];
				if (CVA6Cfg[16543])
					// Trace: core/issue_read_operands.sv:540:9
					tinst_n[i * 32+:32] = issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 0) : (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 3) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 0) : (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 3)) : ((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 0) : (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 3) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 0) : (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 3))) + 31)-:32];
				if (forward_rs1[i])
					// Trace: core/issue_read_operands.sv:545:9
					fu_data_n[(i * ((((12 + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[16503-:32])) + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1))))-:((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1)))) >= (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] + 0))) ? ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1)))) - (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] + 0)))) + 1 : ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] + 0))) - (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1))))) + 1)] = rs1_i[i * CVA6Cfg[17102-:32]+:CVA6Cfg[17102-:32]];
				if (forward_rs2[i])
					// Trace: core/issue_read_operands.sv:548:9
					fu_data_n[(i * ((((12 + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[16503-:32])) + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1)))-:((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1))) >= (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] + 0)) ? ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1))) - (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] + 0))) + 1 : ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] + 0)) - (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1)))) + 1)] = rs2_i[i * CVA6Cfg[17102-:32]+:CVA6Cfg[17102-:32]];
				if ((CVA6Cfg[16471] || (CVA6Cfg[16539] && (OPERANDS_PER_INSTR == 3))) && forward_rs3[i])
					// Trace: core/issue_read_operands.sv:551:9
					fu_data_n[(i * ((((12 + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[16503-:32])) + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1))-:((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1)) >= (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] + 0) ? ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1)) - (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] + 0)) + 1 : ((fu_data_t_fu_data_t_CVA6Cfg[16503-:32] + 0) - (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1))) + 1)] = imm_forward_rs3;
				if (issue_instr_i[(i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 1 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (1 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))])
					// Trace: core/issue_read_operands.sv:556:9
					fu_data_n[(i * ((((12 + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[16503-:32])) + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1))))-:((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1)))) >= (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] + 0))) ? ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1)))) - (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] + 0)))) + 1 : ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] + 0))) - (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1))))) + 1)] = {{CVA6Cfg[17102-:32] - CVA6Cfg[17070-:32] {issue_instr_i[(i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] - 1) - (CVA6Cfg[17070-:32] - 1)) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] - 1) - (CVA6Cfg[17070-:32] - 1))))]}}, issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))))) + ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))))) + 1)) - 1)-:((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))))) + 1)]};
				if (issue_instr_i[(i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 2 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (2 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))])
					// Trace: core/issue_read_operands.sv:564:9
					fu_data_n[(i * ((((12 + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[16503-:32])) + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1))))-:((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1)))) >= (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] + 0))) ? ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1)))) - (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] + 0)))) + 1 : ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] + 0))) - (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1))))) + 1)] = {{CVA6Cfg[17102-:32] - 5 {1'b0}}, issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? 15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? 15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? 15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? 15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1))) + ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)]};
				if ((((issue_instr_i[(i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 3 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (3 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))] && (issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] != 4'd2)) && (issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] != 4'd4)) && (issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] != 4'd10)) && !(CVA6Cfg[16471] && ariane_pkg_is_rs2_fpr(issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)])))
					// Trace: core/issue_read_operands.sv:571:9
					fu_data_n[(i * ((((12 + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[17102-:32]) + fu_data_t_fu_data_t_CVA6Cfg[16503-:32])) + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1)))-:((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1))) >= (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] + 0)) ? ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1))) - (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] + 0))) + 1 : ((fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] + 0)) - (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[17102-:32] + (fu_data_t_fu_data_t_CVA6Cfg[16503-:32] - 1)))) + 1)] = issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) >= (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) + 1 : ((4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + 1)) - 1)-:((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) >= (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) + 1 : ((4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + 1)];
			end
		end
	endgenerate
	// Trace: core/issue_read_operands.sv:578:3
	always @(posedge clk_i or negedge rst_ni)
		// Trace: core/issue_read_operands.sv:579:5
		if (!rst_ni) begin
			// Trace: core/issue_read_operands.sv:580:7
			alu_valid_q <= 1'sb0;
			// Trace: core/issue_read_operands.sv:581:7
			lsu_valid_q <= 1'sb0;
			// Trace: core/issue_read_operands.sv:582:7
			mult_valid_q <= 1'sb0;
			// Trace: core/issue_read_operands.sv:583:7
			fpu_valid_q <= 1'sb0;
			// Trace: core/issue_read_operands.sv:584:7
			fpu_fmt_q <= 1'sb0;
			// Trace: core/issue_read_operands.sv:585:7
			fpu_rm_q <= 1'sb0;
			// Trace: core/issue_read_operands.sv:586:7
			alu2_valid_q <= 1'sb0;
			// Trace: core/issue_read_operands.sv:587:7
			csr_valid_q <= 1'sb0;
			// Trace: core/issue_read_operands.sv:588:7
			branch_valid_q <= 1'sb0;
		end
		else begin
			// Trace: core/issue_read_operands.sv:590:7
			alu_valid_q <= 1'sb0;
			// Trace: core/issue_read_operands.sv:591:7
			lsu_valid_q <= 1'sb0;
			// Trace: core/issue_read_operands.sv:592:7
			mult_valid_q <= 1'sb0;
			// Trace: core/issue_read_operands.sv:593:7
			fpu_valid_q <= 1'sb0;
			// Trace: core/issue_read_operands.sv:594:7
			fpu_fmt_q <= 1'sb0;
			// Trace: core/issue_read_operands.sv:595:7
			fpu_rm_q <= 1'sb0;
			// Trace: core/issue_read_operands.sv:596:7
			alu2_valid_q <= 1'sb0;
			// Trace: core/issue_read_operands.sv:597:7
			csr_valid_q <= 1'sb0;
			// Trace: core/issue_read_operands.sv:598:7
			branch_valid_q <= 1'sb0;
			// Trace: core/issue_read_operands.sv:602:7
			begin : sv2v_autoblock_2
				// Trace: core/issue_read_operands.sv:602:12
				reg [31:0] i;
				// Trace: core/issue_read_operands.sv:602:12
				for (i = 0; i < CVA6Cfg[16841-:32]; i = i + 1)
					begin
						// Trace: core/issue_read_operands.sv:603:9
						if ((!issue_instr_i[(i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) : (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) : (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))] && issue_instr_valid_i[i]) && issue_ack_o[i])
							// Trace: core/issue_read_operands.sv:604:11
							case (issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)])
								4'd3:
									// Trace: core/issue_read_operands.sv:606:15
									if (CVA6Cfg[16874] && !fus_busy[(i * 12) + 7])
										// Trace: core/issue_read_operands.sv:607:17
										alu2_valid_q[i] <= 1'b1;
									else
										// Trace: core/issue_read_operands.sv:609:17
										alu_valid_q[i] <= 1'b1;
								4'd4:
									// Trace: core/issue_read_operands.sv:613:15
									branch_valid_q[i] <= 1'b1;
								4'd5:
									// Trace: core/issue_read_operands.sv:616:15
									mult_valid_q[i] <= 1'b1;
								4'd1, 4'd2:
									// Trace: core/issue_read_operands.sv:619:15
									lsu_valid_q[i] <= 1'b1;
								4'd6:
									// Trace: core/issue_read_operands.sv:622:15
									csr_valid_q[i] <= 1'b1;
								default:
									// Trace: core/issue_read_operands.sv:625:15
									if ((issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] == 4'd7) && CVA6Cfg[16471]) begin
										// Trace: core/issue_read_operands.sv:626:17
										fpu_valid_q[i] <= 1'b1;
										// Trace: core/issue_read_operands.sv:627:17
										fpu_fmt_q <= orig_instr[26-:2];
										// Trace: core/issue_read_operands.sv:628:17
										fpu_rm_q <= orig_instr[14-:3];
									end
									else if ((issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] == 4'd8) && CVA6Cfg[16471]) begin
										// Trace: core/issue_read_operands.sv:630:17
										fpu_valid_q[i] <= 1'b1;
										// Trace: core/issue_read_operands.sv:631:17
										fpu_fmt_q <= orig_instr[13-:2];
										// Trace: core/issue_read_operands.sv:632:17
										fpu_rm_q <= {2'b00, orig_instr[14]};
									end
							endcase
					end
			end
			if (flush_i) begin
				// Trace: core/issue_read_operands.sv:641:9
				alu_valid_q <= 1'sb0;
				// Trace: core/issue_read_operands.sv:642:9
				lsu_valid_q <= 1'sb0;
				// Trace: core/issue_read_operands.sv:643:9
				mult_valid_q <= 1'sb0;
				// Trace: core/issue_read_operands.sv:644:9
				fpu_valid_q <= 1'sb0;
				// Trace: core/issue_read_operands.sv:645:9
				alu2_valid_q <= 1'sb0;
				// Trace: core/issue_read_operands.sv:646:9
				csr_valid_q <= 1'sb0;
				// Trace: core/issue_read_operands.sv:647:9
				branch_valid_q <= 1'sb0;
			end
		end
	// Trace: core/issue_read_operands.sv:652:3
	generate
		if (CVA6Cfg[16539]) begin : genblk6
			// Trace: core/issue_read_operands.sv:653:5
			always @(posedge clk_i or negedge rst_ni)
				// Trace: core/issue_read_operands.sv:654:7
				if (!rst_ni) begin
					// Trace: core/issue_read_operands.sv:655:9
					cvxif_valid_q <= 1'sb0;
					// Trace: core/issue_read_operands.sv:656:9
					cvxif_off_instr_q <= 32'b00000000000000000000000000000000;
				end
				else begin
					// Trace: core/issue_read_operands.sv:658:9
					cvxif_valid_q <= 1'sb0;
					// Trace: core/issue_read_operands.sv:659:9
					cvxif_off_instr_q <= 32'b00000000000000000000000000000000;
					// Trace: core/issue_read_operands.sv:660:9
					begin : sv2v_autoblock_3
						// Trace: core/issue_read_operands.sv:660:14
						reg [31:0] i;
						// Trace: core/issue_read_operands.sv:660:14
						for (i = 0; i < CVA6Cfg[16841-:32]; i = i + 1)
							begin
								// Trace: core/issue_read_operands.sv:661:11
								if ((!issue_instr_i[(i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) : (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) : (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))] && issue_instr_valid_i[i]) && issue_ack_o[i])
									// Trace: core/issue_read_operands.sv:662:13
									case (issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)])
										4'd9: begin
											// Trace: core/issue_read_operands.sv:664:17
											cvxif_valid_q[i] <= 1'b1;
											// Trace: core/issue_read_operands.sv:665:17
											cvxif_off_instr_q <= orig_instr[i];
										end
										default:
											;
									endcase
							end
					end
					if (flush_i) begin
						// Trace: core/issue_read_operands.sv:672:11
						cvxif_valid_q <= 1'sb0;
						// Trace: core/issue_read_operands.sv:673:11
						cvxif_off_instr_q <= 32'b00000000000000000000000000000000;
					end
				end
		end
	endgenerate
	// Trace: core/issue_read_operands.sv:680:3
	always @(*) begin : gen_check_waw_dependencies
		if (_sv2v_0)
			;
		// Trace: core/issue_read_operands.sv:681:5
		stall_waw = 1'sb1;
		// Trace: core/issue_read_operands.sv:682:5
		begin : sv2v_autoblock_4
			// Trace: core/issue_read_operands.sv:682:10
			reg [31:0] i;
			// Trace: core/issue_read_operands.sv:682:10
			for (i = 0; i < CVA6Cfg[16841-:32]; i = i + 1)
				begin
					// Trace: core/issue_read_operands.sv:683:7
					if (issue_instr_valid_i[i] && !fu_busy[i]) begin
						// Trace: core/issue_read_operands.sv:688:9
						if ((CVA6Cfg[16471] && ariane_pkg_is_rd_fpr(issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)]) ? rd_clobber_fpr_i[issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] * 4+:4] == 4'd0 : rd_clobber_gpr_i[issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] * 4+:4] == 4'd0))
							// Trace: core/issue_read_operands.sv:692:11
							stall_waw[i] = 1'b0;
						begin : sv2v_autoblock_5
							// Trace: core/issue_read_operands.sv:696:14
							reg [31:0] c;
							// Trace: core/issue_read_operands.sv:696:14
							for (c = 0; c < CVA6Cfg[16873-:32]; c = c + 1)
								begin
									// Trace: core/issue_read_operands.sv:697:11
									if ((CVA6Cfg[16471] && ariane_pkg_is_rd_fpr(issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)]) ? we_fpr_i[c] && (waddr_i[c * 5+:5] == issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? 5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? 5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? 5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? 5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1))) + ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)]) : we_gpr_i[c] && (waddr_i[c * 5+:5] == issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? 5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? 5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? 5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? 5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1))) + ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)])))
										// Trace: core/issue_read_operands.sv:701:13
										stall_waw[i] = 1'b0;
								end
						end
						if (i > 0) begin
							begin
								// Trace: core/issue_read_operands.sv:705:11
								if ((issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? 5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? 5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? 5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? 5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1))) + ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] == issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((i - 1) * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? 5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? 5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)) : ((((i - 1) * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? 5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? 5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1))) + ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)]) && (issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? 5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? 5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? 5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? 5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1))) + ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (5 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] != {5 {1'sb0}}))
									// Trace: core/issue_read_operands.sv:706:13
									stall_waw[i] = 1'b1;
							end
						end
					end
				end
		end
	end
	// Trace: core/issue_read_operands.sv:715:3
	always @(*) begin : issue_scoreboard
		if (_sv2v_0)
			;
		// Trace: core/issue_read_operands.sv:716:5
		begin : sv2v_autoblock_6
			// Trace: core/issue_read_operands.sv:716:10
			reg [31:0] i;
			// Trace: core/issue_read_operands.sv:716:10
			for (i = 0; i < CVA6Cfg[16841-:32]; i = i + 1)
				begin
					// Trace: core/issue_read_operands.sv:718:7
					issue_ack[i] = 1'b0;
					// Trace: core/issue_read_operands.sv:721:7
					if (issue_instr_valid_i[i] && !fu_busy[i]) begin
						// Trace: core/issue_read_operands.sv:722:9
						if (!stall_raw[i] && !stall_waw[i])
							// Trace: core/issue_read_operands.sv:723:11
							issue_ack[i] = 1'b1;
						if (issue_instr_i[(i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) : (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) : (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))])
							// Trace: core/issue_read_operands.sv:731:11
							issue_ack[i] = 1'b1;
						if (issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] == 4'd0)
							// Trace: core/issue_read_operands.sv:735:11
							issue_ack[i] = 1'b1;
					end
				end
		end
		if (CVA6Cfg[16874]) begin
			begin
				// Trace: core/issue_read_operands.sv:741:7
				if (!issue_ack[0])
					// Trace: core/issue_read_operands.sv:742:9
					issue_ack[1] = 1'b0;
			end
		end
		// Trace: core/issue_read_operands.sv:745:5
		issue_ack_o = issue_ack;
		if ((issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 0 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : ((0 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] == 4'd9) && !(x_transaction_accepted_o || x_transaction_rejected))
			// Trace: core/issue_read_operands.sv:748:7
			issue_ack_o[0] = 1'b0;
	end
	// Trace: core/issue_read_operands.sv:755:3
	wire [(CVA6Cfg[16433-:32] * CVA6Cfg[17102-:32]) - 1:0] rdata;
	// Trace: core/issue_read_operands.sv:756:3
	wire [(CVA6Cfg[16433-:32] * 5) - 1:0] raddr_pack;
	// Trace: core/issue_read_operands.sv:759:3
	wire [(CVA6Cfg[16873-:32] * 5) - 1:0] waddr_pack;
	// Trace: core/issue_read_operands.sv:760:3
	wire [(CVA6Cfg[16873-:32] * CVA6Cfg[17102-:32]) - 1:0] wdata_pack;
	// Trace: core/issue_read_operands.sv:761:3
	wire [CVA6Cfg[16873-:32] - 1:0] we_pack;
	// Trace: core/issue_read_operands.sv:763:3
	genvar _gv_i_37;
	generate
		for (_gv_i_37 = 0; _gv_i_37 < CVA6Cfg[16841-:32]; _gv_i_37 = _gv_i_37 + 1) begin : genblk7
			localparam i = _gv_i_37;
			// Trace: core/issue_read_operands.sv:764:5
			assign raddr_pack[((i * OPERANDS_PER_INSTR) + 0) * 5+:5] = issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? 15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? 15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? 15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? 15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1))) + ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)];
			// Trace: core/issue_read_operands.sv:765:5
			assign raddr_pack[((i * OPERANDS_PER_INSTR) + 1) * 5+:5] = issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? 10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? 10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? 10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? 10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1))) + ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)];
			if (OPERANDS_PER_INSTR == 3) begin : genblk1
				// Trace: core/issue_read_operands.sv:767:7
				assign raddr_pack[((i * OPERANDS_PER_INSTR) + 2) * 5+:5] = issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5) : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) + (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1))) + 1 : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5))) + 1)) - 1) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5) : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) + (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1))) + 1 : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5))) + 1)) - 1)) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5) : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) + (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1))) + 1 : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5))) + 1)) - 1) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5) : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) + (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1))) + 1 : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5))) + 1)) - 1))) + (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1))) + 1 : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5))) + 1)) - 1)-:(((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1))) + 1 : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5))) + 1)];
			end
		end
	endgenerate
	// Trace: core/issue_read_operands.sv:771:3
	genvar _gv_i_38;
	generate
		for (_gv_i_38 = 0; _gv_i_38 < CVA6Cfg[16873-:32]; _gv_i_38 = _gv_i_38 + 1) begin : gen_write_back_port
			localparam i = _gv_i_38;
			// Trace: core/issue_read_operands.sv:772:5
			assign waddr_pack[i * 5+:5] = waddr_i[i * 5+:5];
			// Trace: core/issue_read_operands.sv:773:5
			assign wdata_pack[i * CVA6Cfg[17102-:32]+:CVA6Cfg[17102-:32]] = wdata_i[i * CVA6Cfg[17102-:32]+:CVA6Cfg[17102-:32]];
			// Trace: core/issue_read_operands.sv:774:5
			assign we_pack[i] = we_gpr_i[i];
		end
	endgenerate
	// Trace: core/issue_read_operands.sv:776:3
	generate
		if (CVA6Cfg[16876]) begin : gen_fpga_regfile
			// Trace: core/issue_read_operands.sv:777:5
			ariane_regfile_fpga #(
				.CVA6Cfg(CVA6Cfg),
				.DATA_WIDTH(CVA6Cfg[17102-:32]),
				.NR_READ_PORTS(CVA6Cfg[16433-:32]),
				.ZERO_REG_ZERO(1)
			) i_ariane_regfile_fpga(
				.test_en_i(1'b0),
				.raddr_i(raddr_pack),
				.rdata_o(rdata),
				.waddr_i(waddr_pack),
				.wdata_i(wdata_pack),
				.we_i(we_pack),
				.clk_i(clk_i),
				.rst_ni(rst_ni)
			);
		end
		else begin : gen_asic_regfile
			// Trace: core/issue_read_operands.sv:792:5
			ariane_regfile #(
				.CVA6Cfg(CVA6Cfg),
				.DATA_WIDTH(CVA6Cfg[17102-:32]),
				.NR_READ_PORTS(CVA6Cfg[16433-:32]),
				.ZERO_REG_ZERO(1)
			) i_ariane_regfile(
				.test_en_i(1'b0),
				.raddr_i(raddr_pack),
				.rdata_o(rdata),
				.waddr_i(waddr_pack),
				.wdata_i(wdata_pack),
				.we_i(we_pack),
				.clk_i(clk_i),
				.rst_ni(rst_ni)
			);
		end
	endgenerate
	// Trace: core/issue_read_operands.sv:811:3
	wire [(3 * CVA6Cfg[16469-:32]) - 1:0] fprdata;
	// Trace: core/issue_read_operands.sv:814:3
	reg [14:0] fp_raddr_pack;
	// Trace: core/issue_read_operands.sv:815:3
	wire [(CVA6Cfg[16873-:32] * CVA6Cfg[17102-:32]) - 1:0] fp_wdata_pack;
	// Trace: core/issue_read_operands.sv:817:3
	always @(*) begin : assign_fp_raddr_pack
		if (_sv2v_0)
			;
		// Trace: core/issue_read_operands.sv:818:5
		fp_raddr_pack = {issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 0 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5) : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) + (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1))) + 1 : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5))) + 1)) - 1) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5) : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) + (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1))) + 1 : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5))) + 1)) - 1)) : ((0 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5) : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) + (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1))) + 1 : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5))) + 1)) - 1) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5) : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) + (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1))) + 1 : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5))) + 1)) - 1))) + (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1))) + 1 : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5))) + 1)) - 1)-:(((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1))) + 1 : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5))) + 1)], issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 0 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? 10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? 10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)) : ((0 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? 10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? 10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1))) + ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)], issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 0 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? 15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? 15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)) : ((0 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? 15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? 15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1))) + ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)]};
		// Trace: core/issue_read_operands.sv:822:5
		if (CVA6Cfg[16874]) begin
			begin
				// Trace: core/issue_read_operands.sv:823:7
				if (!(|{issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 0 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : ((0 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] == 4'd7, issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 0 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : ((0 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] == 4'd8}))
					// Trace: core/issue_read_operands.sv:824:9
					fp_raddr_pack = {issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5) : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) + (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1))) + 1 : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5))) + 1)) - 1) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5) : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) + (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1))) + 1 : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5))) + 1)) - 1)) : ((((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5) : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) + (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1))) + 1 : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5))) + 1)) - 1) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5) : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) + (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1))) + 1 : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5))) + 1)) - 1))) + (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1))) + 1 : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5))) + 1)) - 1)-:(((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) >= ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) ? (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1))) + 1 : (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 1)) - ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] - 5))) + 1)], issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? 10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? 10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)) : ((((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? 10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? 10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1))) + ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (10 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)], issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? 15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? 15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)) : ((((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? 15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? 15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) + ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1))) + ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) ? ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4)) + 1 : (((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - 4) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)]};
			end
		end
	end
	// Trace: core/issue_read_operands.sv:831:3
	function automatic [CVA6Cfg[16469-:32] - 1:0] sv2v_cast_76E70;
		input reg [CVA6Cfg[16469-:32] - 1:0] inp;
		sv2v_cast_76E70 = inp;
	endfunction
	generate
		if (CVA6Cfg[16471]) begin : float_regfile_gen
			genvar _gv_i_39;
			for (_gv_i_39 = 0; _gv_i_39 < CVA6Cfg[16873-:32]; _gv_i_39 = _gv_i_39 + 1) begin : gen_fp_wdata_pack
				localparam i = _gv_i_39;
				// Trace: core/issue_read_operands.sv:834:9
				assign fp_wdata_pack[i * CVA6Cfg[17102-:32]+:CVA6Cfg[17102-:32]] = {wdata_i[(i * CVA6Cfg[17102-:32]) + (CVA6Cfg[16469-:32] - 1)-:CVA6Cfg[16469-:32]]};
			end
			if (CVA6Cfg[16876]) begin : gen_fpga_fp_regfile
				// Trace: core/issue_read_operands.sv:837:9
				ariane_regfile_fpga #(
					.CVA6Cfg(CVA6Cfg),
					.DATA_WIDTH(CVA6Cfg[16469-:32]),
					.NR_READ_PORTS(3),
					.ZERO_REG_ZERO(0)
				) i_ariane_fp_regfile_fpga(
					.test_en_i(1'b0),
					.raddr_i(fp_raddr_pack),
					.rdata_o(fprdata),
					.waddr_i(waddr_pack),
					.wdata_i(fp_wdata_pack),
					.we_i(we_fpr_i),
					.clk_i(clk_i),
					.rst_ni(rst_ni)
				);
			end
			else begin : gen_asic_fp_regfile
				// Trace: core/issue_read_operands.sv:852:9
				ariane_regfile #(
					.CVA6Cfg(CVA6Cfg),
					.DATA_WIDTH(CVA6Cfg[16469-:32]),
					.NR_READ_PORTS(3),
					.ZERO_REG_ZERO(0)
				) i_ariane_fp_regfile(
					.test_en_i(1'b0),
					.raddr_i(fp_raddr_pack),
					.rdata_o(fprdata),
					.waddr_i(waddr_pack),
					.wdata_i(fp_wdata_pack),
					.we_i(we_fpr_i),
					.clk_i(clk_i),
					.rst_ni(rst_ni)
				);
			end
		end
		else begin : no_fpr_gen
			// Trace: core/issue_read_operands.sv:868:7
			assign fprdata = {3 {sv2v_cast_76E70(1'sb0)}};
		end
	endgenerate
	// Trace: core/issue_read_operands.sv:872:3
	generate
		if (OPERANDS_PER_INSTR == 3) begin : gen_operand_c
			// Trace: core/issue_read_operands.sv:873:5
			assign operand_c_fpr = {{CVA6Cfg[17102-:32] - CVA6Cfg[16469-:32] {1'b0}}, fprdata[2 * CVA6Cfg[16469-:32]+:CVA6Cfg[16469-:32]]};
		end
		else begin : genblk11
			// Trace: core/issue_read_operands.sv:875:5
			assign operand_c_fpr = fprdata[2 * CVA6Cfg[16469-:32]+:CVA6Cfg[16469-:32]];
		end
	endgenerate
	// Trace: core/issue_read_operands.sv:878:3
	genvar _gv_i_40;
	generate
		for (_gv_i_40 = 0; _gv_i_40 < CVA6Cfg[16841-:32]; _gv_i_40 = _gv_i_40 + 1) begin : genblk12
			localparam i = _gv_i_40;
			if (OPERANDS_PER_INSTR == 3) begin : gen_operand_c
				// Trace: core/issue_read_operands.sv:880:7
				assign operand_c_gpr[i * (rs3_len_t_CVA6Cfg[16433-:32] == 3 ? rs3_len_t_CVA6Cfg[17102-:32] : rs3_len_t_CVA6Cfg[16469-:32])+:(rs3_len_t_CVA6Cfg[16433-:32] == 3 ? rs3_len_t_CVA6Cfg[17102-:32] : rs3_len_t_CVA6Cfg[16469-:32])] = rdata[((i * OPERANDS_PER_INSTR) + 2) * CVA6Cfg[17102-:32]+:CVA6Cfg[17102-:32]];
			end
			// Trace: core/issue_read_operands.sv:883:5
			assign operand_a_regfile[i * CVA6Cfg[17102-:32]+:CVA6Cfg[17102-:32]] = (CVA6Cfg[16471] && ariane_pkg_is_rs1_fpr(issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)]) ? {{CVA6Cfg[17102-:32] - CVA6Cfg[16469-:32] {1'b0}}, fprdata[0+:CVA6Cfg[16469-:32]]} : rdata[((i * OPERANDS_PER_INSTR) + 0) * CVA6Cfg[17102-:32]+:CVA6Cfg[17102-:32]]);
			// Trace: core/issue_read_operands.sv:886:5
			assign operand_b_regfile[i * CVA6Cfg[17102-:32]+:CVA6Cfg[17102-:32]] = (CVA6Cfg[16471] && ariane_pkg_is_rs2_fpr(issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)]) ? {{CVA6Cfg[17102-:32] - CVA6Cfg[16469-:32] {1'b0}}, fprdata[CVA6Cfg[16469-:32]+:CVA6Cfg[16469-:32]]} : rdata[((i * OPERANDS_PER_INSTR) + 1) * CVA6Cfg[17102-:32]+:CVA6Cfg[17102-:32]]);
			// Trace: core/issue_read_operands.sv:889:5
			assign operand_c_regfile[i * (rs3_len_t_CVA6Cfg[16433-:32] == 3 ? rs3_len_t_CVA6Cfg[17102-:32] : rs3_len_t_CVA6Cfg[16469-:32])+:(rs3_len_t_CVA6Cfg[16433-:32] == 3 ? rs3_len_t_CVA6Cfg[17102-:32] : rs3_len_t_CVA6Cfg[16469-:32])] = (OPERANDS_PER_INSTR == 3 ? (CVA6Cfg[16471] && ariane_pkg_is_imm_fpr(issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((i * ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4))) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((15 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)]) ? operand_c_fpr : operand_c_gpr[i * (rs3_len_t_CVA6Cfg[16433-:32] == 3 ? rs3_len_t_CVA6Cfg[17102-:32] : rs3_len_t_CVA6Cfg[16469-:32])+:(rs3_len_t_CVA6Cfg[16433-:32] == 3 ? rs3_len_t_CVA6Cfg[17102-:32] : rs3_len_t_CVA6Cfg[16469-:32])]) : operand_c_fpr);
		end
	endgenerate
	// Trace: core/issue_read_operands.sv:897:3
	// removed localparam type ariane_pkg_cf_t
	always @(posedge clk_i or negedge rst_ni)
		// Trace: core/issue_read_operands.sv:898:5
		if (!rst_ni) begin
			// Trace: core/issue_read_operands.sv:899:7
			fu_data_q <= 1'sb0;
			// Trace: core/issue_read_operands.sv:900:7
			if (CVA6Cfg[16543])
				// Trace: core/issue_read_operands.sv:901:9
				tinst_q <= 1'sb0;
			// Trace: core/issue_read_operands.sv:903:7
			pc_o <= 1'sb0;
			// Trace: core/issue_read_operands.sv:904:7
			is_compressed_instr_o <= 1'b0;
			// Trace: core/issue_read_operands.sv:905:7
			branch_predict_o <= {3'd0, {CVA6Cfg[17070-:32] {1'b0}}};
			// Trace: core/issue_read_operands.sv:906:7
			x_transaction_rejected_o <= 1'b0;
		end
		else begin
			// Trace: core/issue_read_operands.sv:908:7
			fu_data_q <= fu_data_n;
			// Trace: core/issue_read_operands.sv:909:7
			if (CVA6Cfg[16543])
				// Trace: core/issue_read_operands.sv:910:9
				tinst_q <= tinst_n;
			if (CVA6Cfg[16874]) begin
				begin
					// Trace: core/issue_read_operands.sv:913:9
					if (issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : ((((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] == 4'd4) begin
						// Trace: core/issue_read_operands.sv:914:11
						pc_o <= issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))))) : ((((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))))) + ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))))) + 1)) - 1)-:((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))))) + 1)];
						// Trace: core/issue_read_operands.sv:915:11
						is_compressed_instr_o <= issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 4 : ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 0)];
						// Trace: core/issue_read_operands.sv:916:11
						branch_predict_o <= issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4 : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) : ((((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 5 : 1 - (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4)) + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4 : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))) + (((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4) >= 5 ? (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 0 : 6 - ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))) - 1)-:(((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4) >= 5 ? (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 0 : 6 - ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))];
					end
				end
			end
			if (issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 0 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : ((0 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] == 4'd4) begin
				// Trace: core/issue_read_operands.sv:920:9
				pc_o <= issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 0 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))))) : ((0 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))))) + ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))))) + 1)) - 1)-:((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) >= (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))))) + 1 : ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) - (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32] + (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))))) + 1)];
				// Trace: core/issue_read_operands.sv:921:9
				is_compressed_instr_o <= issue_instr_i[0 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 4 : ((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 0)];
				// Trace: core/issue_read_operands.sv:922:9
				branch_predict_o <= issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 0 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4 : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)) : ((0 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4 : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))) + (((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4) >= 5 ? (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 0 : 6 - ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))) - 1)-:(((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4) >= 5 ? (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 0 : 6 - ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))];
			end
			// Trace: core/issue_read_operands.sv:924:7
			x_transaction_rejected_o <= 1'b0;
			if (issue_instr_i[((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 0 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) : ((0 + ((((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) >= 0 ? 27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))) : (((((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[16503-:32]) + 27) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + 4) + ((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33))) + (3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32])) + 4) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))))) + ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)) - 1)-:((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) >= (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) ? ((27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4))))) - (23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5)))))) + 1 : ((23 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 5))))) - (27 + (scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + (4 + (((((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33) >= 0 ? ((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 34 : 1 - (((scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32] + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17102-:32]) + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17006-:32]) + 33)) + ((3 + scoreboard_entry_t_scoreboard_entry_t_CVA6Cfg[17070-:32]) + 4)))))) + 1)] == 4'd9)
				// Trace: core/issue_read_operands.sv:926:9
				x_transaction_rejected_o <= x_transaction_rejected;
		end
	// Trace: core/issue_read_operands.sv:932:3
	// Trace: core/issue_read_operands.sv:949:3
	// Trace: core/issue_read_operands.sv:955:3
	genvar _gv_i_41;
	generate
		for (_gv_i_41 = 0; _gv_i_41 < CVA6Cfg[16841-:32]; _gv_i_41 = _gv_i_41 + 1) begin : genblk13
			localparam i = _gv_i_41;
			// Trace: core/issue_read_operands.sv:956:5
			// removed an assertion item
			// assert property (@(posedge clk_i) 
			// 	(branch_valid_q |-> !$isunknown(fu_data_q[i].operand_a) && !$isunknown(fu_data_q[i].operand_b))
			// ) else begin
			// 	// Trace: core/issue_read_operands.sv:961:10
			// 	$warning("Got unknown value in one of the operands");
			// end
		end
	endgenerate
	initial _sv2v_0 = 0;
endmodule
