module store_buffer_AA2E5_FDA9C (
	clk_i,
	rst_ni,
	flush_i,
	stall_st_pending_i,
	no_st_pending_o,
	store_buffer_empty_o,
	page_offset_i,
	page_offset_matches_o,
	commit_i,
	commit_ready_o,
	ready_o,
	valid_i,
	valid_without_flush_i,
	paddr_i,
	rvfi_mem_paddr_o,
	data_i,
	be_i,
	data_size_i,
	req_port_i,
	req_port_o
);
	// removed localparam type dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg_type
	parameter [17102:0] dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg = 0;
	// removed localparam type dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg_type
	parameter [17102:0] dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg = 0;
	reg _sv2v_0;
	// removed import ariane_pkg::*;
	// Trace: core/store_buffer.sv:20:15
	localparam config_pkg_NrMaxRules = 16;
	// removed localparam type config_pkg_cache_type_t
	// removed localparam type config_pkg_noc_type_e
	// removed localparam type config_pkg_vm_mode_t
	// removed localparam type config_pkg_cva6_cfg_t
	localparam [17102:0] config_pkg_cva6_cfg_empty = 17103'd0;
	parameter [17102:0] CVA6Cfg = config_pkg_cva6_cfg_empty;
	// Trace: core/store_buffer.sv:21:20
	// removed localparam type dcache_req_i_t
	// Trace: core/store_buffer.sv:22:20
	// removed localparam type dcache_req_o_t
	// Trace: core/store_buffer.sv:24:5
	input wire clk_i;
	// Trace: core/store_buffer.sv:25:5
	input wire rst_ni;
	// Trace: core/store_buffer.sv:26:5
	input wire flush_i;
	// Trace: core/store_buffer.sv:28:5
	input wire stall_st_pending_i;
	// Trace: core/store_buffer.sv:29:5
	output reg no_st_pending_o;
	// Trace: core/store_buffer.sv:30:5
	output wire store_buffer_empty_o;
	// Trace: core/store_buffer.sv:32:5
	input wire [11:0] page_offset_i;
	// Trace: core/store_buffer.sv:33:5
	output reg page_offset_matches_o;
	// Trace: core/store_buffer.sv:35:5
	input wire commit_i;
	// Trace: core/store_buffer.sv:36:5
	output reg commit_ready_o;
	// Trace: core/store_buffer.sv:37:5
	output reg ready_o;
	// Trace: core/store_buffer.sv:40:5
	input wire valid_i;
	// Trace: core/store_buffer.sv:41:5
	input wire valid_without_flush_i;
	// Trace: core/store_buffer.sv:43:5
	input wire [CVA6Cfg[17038-:32] - 1:0] paddr_i;
	// Trace: core/store_buffer.sv:44:5
	output wire [CVA6Cfg[17038-:32] - 1:0] rvfi_mem_paddr_o;
	// Trace: core/store_buffer.sv:45:5
	input wire [CVA6Cfg[17102-:32] - 1:0] data_i;
	// Trace: core/store_buffer.sv:46:5
	input wire [(CVA6Cfg[17102-:32] / 8) - 1:0] be_i;
	// Trace: core/store_buffer.sv:47:5
	input wire [1:0] data_size_i;
	// Trace: core/store_buffer.sv:50:5
	input wire [(((2 + dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[1124-:32]) + dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[17102-:32]) + dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[900-:32]) - 1:0] req_port_i;
	// Trace: core/store_buffer.sv:51:5
	output reg [(((((((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1028-:32] + dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[996-:32]) + dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32]) + dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32]) + 2) + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8)) + 2) + dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32]) + 1:0] req_port_o;
	// Trace: core/store_buffer.sv:57:3
	localparam [2:0] ariane_pkg_DEPTH_SPEC = 'd4;
	reg [((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? (ariane_pkg_DEPTH_SPEC * (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 3)) - 1 : (ariane_pkg_DEPTH_SPEC * (1 - (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2))) + (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 1)):((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? 0 : ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2)] speculative_queue_n;
	reg [((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? (ariane_pkg_DEPTH_SPEC * (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 3)) - 1 : (ariane_pkg_DEPTH_SPEC * (1 - (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2))) + (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 1)):((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? 0 : ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2)] speculative_queue_q;
	localparam [2:0] ariane_pkg_DEPTH_COMMIT = 'd4;
	reg [((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? (ariane_pkg_DEPTH_COMMIT * (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 3)) - 1 : (ariane_pkg_DEPTH_COMMIT * (1 - (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2))) + (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 1)):((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? 0 : ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2)] commit_queue_n;
	reg [((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? (ariane_pkg_DEPTH_COMMIT * (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 3)) - 1 : (ariane_pkg_DEPTH_COMMIT * (1 - (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2))) + (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 1)):((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? 0 : ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2)] commit_queue_q;
	// Trace: core/store_buffer.sv:70:3
	reg [$clog2(3'd4):0] speculative_status_cnt_n;
	reg [$clog2(3'd4):0] speculative_status_cnt_q;
	// Trace: core/store_buffer.sv:71:3
	reg [$clog2(3'd4):0] commit_status_cnt_n;
	reg [$clog2(3'd4):0] commit_status_cnt_q;
	// Trace: core/store_buffer.sv:73:3
	reg [$clog2(3'd4) - 1:0] speculative_read_pointer_n;
	reg [$clog2(3'd4) - 1:0] speculative_read_pointer_q;
	// Trace: core/store_buffer.sv:74:3
	reg [$clog2(3'd4) - 1:0] speculative_write_pointer_n;
	reg [$clog2(3'd4) - 1:0] speculative_write_pointer_q;
	// Trace: core/store_buffer.sv:76:3
	reg [$clog2(3'd4) - 1:0] commit_read_pointer_n;
	reg [$clog2(3'd4) - 1:0] commit_read_pointer_q;
	// Trace: core/store_buffer.sv:77:3
	reg [$clog2(3'd4) - 1:0] commit_write_pointer_n;
	reg [$clog2(3'd4) - 1:0] commit_write_pointer_q;
	// Trace: core/store_buffer.sv:79:3
	assign store_buffer_empty_o = (speculative_status_cnt_q == 0) & no_st_pending_o;
	// Trace: core/store_buffer.sv:83:3
	always @(*) begin : core_if
		// Trace: core/store_buffer.sv:84:5
		reg [$clog2(3'd4):0] speculative_status_cnt;
		if (_sv2v_0)
			;
		// Trace: core/store_buffer.sv:85:5
		speculative_status_cnt = speculative_status_cnt_q;
		// Trace: core/store_buffer.sv:88:5
		speculative_status_cnt_n = speculative_status_cnt_q;
		// Trace: core/store_buffer.sv:89:5
		speculative_read_pointer_n = speculative_read_pointer_q;
		// Trace: core/store_buffer.sv:90:5
		speculative_write_pointer_n = speculative_write_pointer_q;
		// Trace: core/store_buffer.sv:91:5
		speculative_queue_n = speculative_queue_q;
		// Trace: core/store_buffer.sv:94:5
		if (valid_i) begin
			// Trace: core/store_buffer.sv:95:7
			speculative_queue_n[((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? (speculative_write_pointer_q * ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 3 : 1 - (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2))) + ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2)) : (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) - (CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2)))) : (((speculative_write_pointer_q * ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 3 : 1 - (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2))) + ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2)) : (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) - (CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))))) + ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) >= (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 3)) ? ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 3))) + 1 : ((CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 3)) - (CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2)))) + 1)) - 1)-:((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) >= (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 3)) ? ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 3))) + 1 : ((CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 3)) - (CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2)))) + 1)] = paddr_i;
			// Trace: core/store_buffer.sv:96:7
			speculative_queue_n[((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? (speculative_write_pointer_q * ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 3 : 1 - (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2))) + ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2) : (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) - (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) : (((speculative_write_pointer_q * ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 3 : 1 - (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2))) + ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2) : (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) - (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2)))) + ((CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2)) >= ((CVA6Cfg[17102-:32] / 8) + 3) ? ((CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2)) - ((CVA6Cfg[17102-:32] / 8) + 3)) + 1 : (((CVA6Cfg[17102-:32] / 8) + 3) - (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) + 1)) - 1)-:((CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2)) >= ((CVA6Cfg[17102-:32] / 8) + 3) ? ((CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2)) - ((CVA6Cfg[17102-:32] / 8) + 3)) + 1 : (((CVA6Cfg[17102-:32] / 8) + 3) - (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) + 1)] = data_i;
			// Trace: core/store_buffer.sv:97:7
			speculative_queue_n[((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? (speculative_write_pointer_q * ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 3 : 1 - (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2))) + ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? (CVA6Cfg[17102-:32] / 8) + 2 : (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) - ((CVA6Cfg[17102-:32] / 8) + 2)) : (((speculative_write_pointer_q * ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 3 : 1 - (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2))) + ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? (CVA6Cfg[17102-:32] / 8) + 2 : (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) - ((CVA6Cfg[17102-:32] / 8) + 2))) + (((CVA6Cfg[17102-:32] / 8) + 2) >= 3 ? (CVA6Cfg[17102-:32] / 8) + 0 : 4 - ((CVA6Cfg[17102-:32] / 8) + 2))) - 1)-:(((CVA6Cfg[17102-:32] / 8) + 2) >= 3 ? (CVA6Cfg[17102-:32] / 8) + 0 : 4 - ((CVA6Cfg[17102-:32] / 8) + 2))] = be_i;
			// Trace: core/store_buffer.sv:98:7
			speculative_queue_n[((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? (speculative_write_pointer_q * ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 3 : 1 - (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2))) + ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? 2 : ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 0) : ((speculative_write_pointer_q * ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 3 : 1 - (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2))) + ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? 2 : ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 0)) + 1)-:2] = data_size_i;
			// Trace: core/store_buffer.sv:99:7
			speculative_queue_n[(speculative_write_pointer_q * ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 3 : 1 - (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2))) + ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? 0 : ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2)] = 1'b1;
			// Trace: core/store_buffer.sv:101:7
			speculative_write_pointer_n = speculative_write_pointer_q + 1'b1;
			// Trace: core/store_buffer.sv:102:7
			speculative_status_cnt = speculative_status_cnt + 1;
		end
		if (commit_i) begin
			// Trace: core/store_buffer.sv:109:7
			speculative_queue_n[(speculative_read_pointer_q * ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 3 : 1 - (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2))) + ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? 0 : ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2)] = 1'b0;
			// Trace: core/store_buffer.sv:111:7
			speculative_read_pointer_n = speculative_read_pointer_q + 1'b1;
			// Trace: core/store_buffer.sv:112:7
			speculative_status_cnt = speculative_status_cnt - 1;
		end
		// Trace: core/store_buffer.sv:115:5
		speculative_status_cnt_n = speculative_status_cnt;
		if (flush_i) begin
			// Trace: core/store_buffer.sv:120:7
			begin : sv2v_autoblock_1
				// Trace: core/store_buffer.sv:120:12
				reg [31:0] i;
				// Trace: core/store_buffer.sv:120:12
				for (i = 0; i < ariane_pkg_DEPTH_SPEC; i = i + 1)
					begin
						// Trace: core/store_buffer.sv:120:53
						speculative_queue_n[(i * ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 3 : 1 - (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2))) + ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? 0 : ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2)] = 1'b0;
					end
			end
			// Trace: core/store_buffer.sv:122:7
			speculative_write_pointer_n = speculative_read_pointer_q;
			// Trace: core/store_buffer.sv:124:7
			speculative_status_cnt_n = 'b0;
		end
		// Trace: core/store_buffer.sv:128:5
		ready_o = (speculative_status_cnt_n < ariane_pkg_DEPTH_SPEC) || commit_i;
	end
	// Trace: core/store_buffer.sv:137:3
	wire [1:1] sv2v_tmp_DD30F;
	assign sv2v_tmp_DD30F = 1'b0;
	always @(*) req_port_o[1] = sv2v_tmp_DD30F;
	// Trace: core/store_buffer.sv:138:3
	wire [1:1] sv2v_tmp_FEE84;
	assign sv2v_tmp_FEE84 = 1'b1;
	always @(*) req_port_o[1 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1)))] = sv2v_tmp_FEE84;
	// Trace: core/store_buffer.sv:139:3
	wire [1:1] sv2v_tmp_7ADAE;
	assign sv2v_tmp_7ADAE = 1'b0;
	always @(*) req_port_o[0] = sv2v_tmp_7ADAE;
	// Trace: core/store_buffer.sv:142:3
	wire [((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1) >= 2 ? dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 0 : 3 - (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1)) * 1:1] sv2v_tmp_C77FB;
	assign sv2v_tmp_C77FB = 1'sb0;
	always @(*) req_port_o[dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1-:((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1) >= 2 ? dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 0 : 3 - (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1))] = sv2v_tmp_C77FB;
	// Trace: core/store_buffer.sv:144:3
	wire [((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1028-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[996-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1)))))))) >= (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[996-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2))))))) ? ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1028-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[996-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1)))))))) - (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[996-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2)))))))) + 1 : ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[996-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2))))))) - (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1028-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[996-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1))))))))) + 1) * 1:1] sv2v_tmp_FF939;
	assign sv2v_tmp_FF939 = commit_queue_q[((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? (commit_read_pointer_q * ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 3 : 1 - (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2))) + ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - (CVA6Cfg[1028-:32] - 1))) >= ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 1)) ? (CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - (CVA6Cfg[1028-:32] - 1)) : (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - (CVA6Cfg[1028-:32] - 1))) + (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - (CVA6Cfg[1028-:32] - 1))) >= ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 1)) ? (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - (CVA6Cfg[1028-:32] - 1))) - ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 1))) + 1 : (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 1)) - ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - (CVA6Cfg[1028-:32] - 1)))) + 1)) - 1) : (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) - (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - (CVA6Cfg[1028-:32] - 1))) >= ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 1)) ? (CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - (CVA6Cfg[1028-:32] - 1)) : (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - (CVA6Cfg[1028-:32] - 1))) + (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - (CVA6Cfg[1028-:32] - 1))) >= ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 1)) ? (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - (CVA6Cfg[1028-:32] - 1))) - ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 1))) + 1 : (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 1)) - ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - (CVA6Cfg[1028-:32] - 1)))) + 1)) - 1)) : (((commit_read_pointer_q * ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 3 : 1 - (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2))) + ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - (CVA6Cfg[1028-:32] - 1))) >= ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 1)) ? (CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - (CVA6Cfg[1028-:32] - 1)) : (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - (CVA6Cfg[1028-:32] - 1))) + (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - (CVA6Cfg[1028-:32] - 1))) >= ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 1)) ? (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - (CVA6Cfg[1028-:32] - 1))) - ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 1))) + 1 : (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 1)) - ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - (CVA6Cfg[1028-:32] - 1)))) + 1)) - 1) : (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) - (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - (CVA6Cfg[1028-:32] - 1))) >= ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 1)) ? (CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - (CVA6Cfg[1028-:32] - 1)) : (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - (CVA6Cfg[1028-:32] - 1))) + (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - (CVA6Cfg[1028-:32] - 1))) >= ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 1)) ? (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - (CVA6Cfg[1028-:32] - 1))) - ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 1))) + 1 : (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 1)) - ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - (CVA6Cfg[1028-:32] - 1)))) + 1)) - 1))) + (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - (CVA6Cfg[1028-:32] - 1))) >= ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 1)) ? (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - (CVA6Cfg[1028-:32] - 1))) - ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 1))) + 1 : (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 1)) - ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - (CVA6Cfg[1028-:32] - 1)))) + 1)) - 1)-:(((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - (CVA6Cfg[1028-:32] - 1))) >= ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 1)) ? (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - (CVA6Cfg[1028-:32] - 1))) - ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 1))) + 1 : (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 1)) - ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - (CVA6Cfg[1028-:32] - 1)))) + 1)];
	always @(*) req_port_o[dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1028-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[996-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1)))))))-:((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1028-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[996-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1)))))))) >= (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[996-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2))))))) ? ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1028-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[996-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1)))))))) - (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[996-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2)))))))) + 1 : ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[996-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2))))))) - (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1028-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[996-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1))))))))) + 1)] = sv2v_tmp_FF939;
	// Trace: core/store_buffer.sv:146:3
	wire [((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[996-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1))))))) >= (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2)))))) ? ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[996-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1))))))) - (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2))))))) + 1 : ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2)))))) - (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[996-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1)))))))) + 1) * 1:1] sv2v_tmp_32EA6;
	assign sv2v_tmp_32EA6 = commit_queue_q[((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? (commit_read_pointer_q * ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 3 : 1 - (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2))) + ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - ((CVA6Cfg[996-:32] + CVA6Cfg[1028-:32]) - 1))) >= ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - CVA6Cfg[1028-:32])) ? (CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - ((CVA6Cfg[996-:32] + CVA6Cfg[1028-:32]) - 1)) : (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - ((CVA6Cfg[996-:32] + CVA6Cfg[1028-:32]) - 1))) + (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - ((CVA6Cfg[996-:32] + CVA6Cfg[1028-:32]) - 1))) >= ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - CVA6Cfg[1028-:32])) ? (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - ((CVA6Cfg[996-:32] + CVA6Cfg[1028-:32]) - 1))) - ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - CVA6Cfg[1028-:32]))) + 1 : (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - CVA6Cfg[1028-:32])) - ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - ((CVA6Cfg[996-:32] + CVA6Cfg[1028-:32]) - 1)))) + 1)) - 1) : (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) - (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - ((CVA6Cfg[996-:32] + CVA6Cfg[1028-:32]) - 1))) >= ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - CVA6Cfg[1028-:32])) ? (CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - ((CVA6Cfg[996-:32] + CVA6Cfg[1028-:32]) - 1)) : (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - ((CVA6Cfg[996-:32] + CVA6Cfg[1028-:32]) - 1))) + (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - ((CVA6Cfg[996-:32] + CVA6Cfg[1028-:32]) - 1))) >= ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - CVA6Cfg[1028-:32])) ? (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - ((CVA6Cfg[996-:32] + CVA6Cfg[1028-:32]) - 1))) - ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - CVA6Cfg[1028-:32]))) + 1 : (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - CVA6Cfg[1028-:32])) - ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - ((CVA6Cfg[996-:32] + CVA6Cfg[1028-:32]) - 1)))) + 1)) - 1)) : (((commit_read_pointer_q * ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 3 : 1 - (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2))) + ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - ((CVA6Cfg[996-:32] + CVA6Cfg[1028-:32]) - 1))) >= ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - CVA6Cfg[1028-:32])) ? (CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - ((CVA6Cfg[996-:32] + CVA6Cfg[1028-:32]) - 1)) : (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - ((CVA6Cfg[996-:32] + CVA6Cfg[1028-:32]) - 1))) + (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - ((CVA6Cfg[996-:32] + CVA6Cfg[1028-:32]) - 1))) >= ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - CVA6Cfg[1028-:32])) ? (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - ((CVA6Cfg[996-:32] + CVA6Cfg[1028-:32]) - 1))) - ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - CVA6Cfg[1028-:32]))) + 1 : (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - CVA6Cfg[1028-:32])) - ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - ((CVA6Cfg[996-:32] + CVA6Cfg[1028-:32]) - 1)))) + 1)) - 1) : (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) - (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - ((CVA6Cfg[996-:32] + CVA6Cfg[1028-:32]) - 1))) >= ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - CVA6Cfg[1028-:32])) ? (CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - ((CVA6Cfg[996-:32] + CVA6Cfg[1028-:32]) - 1)) : (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - ((CVA6Cfg[996-:32] + CVA6Cfg[1028-:32]) - 1))) + (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - ((CVA6Cfg[996-:32] + CVA6Cfg[1028-:32]) - 1))) >= ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - CVA6Cfg[1028-:32])) ? (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - ((CVA6Cfg[996-:32] + CVA6Cfg[1028-:32]) - 1))) - ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - CVA6Cfg[1028-:32]))) + 1 : (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - CVA6Cfg[1028-:32])) - ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - ((CVA6Cfg[996-:32] + CVA6Cfg[1028-:32]) - 1)))) + 1)) - 1))) + (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - ((CVA6Cfg[996-:32] + CVA6Cfg[1028-:32]) - 1))) >= ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - CVA6Cfg[1028-:32])) ? (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - ((CVA6Cfg[996-:32] + CVA6Cfg[1028-:32]) - 1))) - ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - CVA6Cfg[1028-:32]))) + 1 : (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - CVA6Cfg[1028-:32])) - ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - ((CVA6Cfg[996-:32] + CVA6Cfg[1028-:32]) - 1)))) + 1)) - 1)-:(((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - ((CVA6Cfg[996-:32] + CVA6Cfg[1028-:32]) - 1))) >= ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - CVA6Cfg[1028-:32])) ? (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - ((CVA6Cfg[996-:32] + CVA6Cfg[1028-:32]) - 1))) - ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - CVA6Cfg[1028-:32]))) + 1 : (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - CVA6Cfg[1028-:32])) - ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - ((CVA6Cfg[17038-:32] - 1) - ((CVA6Cfg[996-:32] + CVA6Cfg[1028-:32]) - 1)))) + 1)];
	always @(*) req_port_o[dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[996-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1))))))-:((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[996-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1))))))) >= (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2)))))) ? ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[996-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1))))))) - (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2))))))) + 1 : ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2)))))) - (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[996-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1)))))))) + 1)] = sv2v_tmp_32EA6;
	// Trace: core/store_buffer.sv:149:3
	wire [((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1)))))) >= (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2))))) ? ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1)))))) - (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2)))))) + 1 : ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2))))) - (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1))))))) + 1) * 1:1] sv2v_tmp_29594;
	assign sv2v_tmp_29594 = commit_queue_q[((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? (commit_read_pointer_q * ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 3 : 1 - (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2))) + ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2) : (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) - (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) : (((commit_read_pointer_q * ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 3 : 1 - (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2))) + ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2) : (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) - (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2)))) + ((CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2)) >= ((CVA6Cfg[17102-:32] / 8) + 3) ? ((CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2)) - ((CVA6Cfg[17102-:32] / 8) + 3)) + 1 : (((CVA6Cfg[17102-:32] / 8) + 3) - (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) + 1)) - 1)-:((CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2)) >= ((CVA6Cfg[17102-:32] / 8) + 3) ? ((CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2)) - ((CVA6Cfg[17102-:32] / 8) + 3)) + 1 : (((CVA6Cfg[17102-:32] / 8) + 3) - (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) + 1)];
	always @(*) req_port_o[dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1)))))-:((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1)))))) >= (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2))))) ? ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1)))))) - (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2)))))) + 1 : ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2))))) - (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[900-:32] + (2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1))))))) + 1)] = sv2v_tmp_29594;
	// Trace: core/store_buffer.sv:150:3
	wire [(((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1))) >= (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2)) ? (((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1))) - (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2))) + 1 : ((2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2)) - ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1)))) + 1) * 1:1] sv2v_tmp_C5836;
	assign sv2v_tmp_C5836 = commit_queue_q[((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? (commit_read_pointer_q * ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 3 : 1 - (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2))) + ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? (CVA6Cfg[17102-:32] / 8) + 2 : (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) - ((CVA6Cfg[17102-:32] / 8) + 2)) : (((commit_read_pointer_q * ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 3 : 1 - (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2))) + ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? (CVA6Cfg[17102-:32] / 8) + 2 : (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) - ((CVA6Cfg[17102-:32] / 8) + 2))) + (((CVA6Cfg[17102-:32] / 8) + 2) >= 3 ? (CVA6Cfg[17102-:32] / 8) + 0 : 4 - ((CVA6Cfg[17102-:32] / 8) + 2))) - 1)-:(((CVA6Cfg[17102-:32] / 8) + 2) >= 3 ? (CVA6Cfg[17102-:32] / 8) + 0 : 4 - ((CVA6Cfg[17102-:32] / 8) + 2))];
	always @(*) req_port_o[(dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1))-:(((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1))) >= (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2)) ? (((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1))) - (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2))) + 1 : ((2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2)) - ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1)))) + 1)] = sv2v_tmp_C5836;
	// Trace: core/store_buffer.sv:151:3
	wire [((2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1)) >= (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2) ? ((2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1)) - (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2)) + 1 : ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2) - (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1))) + 1) * 1:1] sv2v_tmp_15C08;
	assign sv2v_tmp_15C08 = commit_queue_q[((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? (commit_read_pointer_q * ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 3 : 1 - (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2))) + ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? 2 : ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 0) : ((commit_read_pointer_q * ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 3 : 1 - (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2))) + ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? 2 : ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 0)) + 1)-:2];
	always @(*) req_port_o[2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1)-:((2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1)) >= (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2) ? ((2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1)) - (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2)) + 1 : ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 2) - (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1))) + 1)] = sv2v_tmp_15C08;
	// Trace: core/store_buffer.sv:153:3
	assign rvfi_mem_paddr_o = commit_queue_n[((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? (commit_read_pointer_n * ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 3 : 1 - (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2))) + ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2)) : (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) - (CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2)))) : (((commit_read_pointer_n * ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 3 : 1 - (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2))) + ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2)) : (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) - (CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))))) + ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) >= (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 3)) ? ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 3))) + 1 : ((CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 3)) - (CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2)))) + 1)) - 1)-:((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) >= (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 3)) ? ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 3))) + 1 : ((CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 3)) - (CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2)))) + 1)];
	// Trace: core/store_buffer.sv:155:3
	always @(*) begin : store_if
		// Trace: core/store_buffer.sv:156:5
		reg [$clog2(3'd4):0] commit_status_cnt;
		if (_sv2v_0)
			;
		// Trace: core/store_buffer.sv:157:5
		commit_status_cnt = commit_status_cnt_q;
		// Trace: core/store_buffer.sv:159:5
		commit_ready_o = commit_status_cnt_q < ariane_pkg_DEPTH_COMMIT;
		// Trace: core/store_buffer.sv:161:5
		no_st_pending_o = commit_status_cnt_q == 0;
		// Trace: core/store_buffer.sv:163:5
		commit_read_pointer_n = commit_read_pointer_q;
		// Trace: core/store_buffer.sv:164:5
		commit_write_pointer_n = commit_write_pointer_q;
		// Trace: core/store_buffer.sv:166:5
		commit_queue_n = commit_queue_q;
		// Trace: core/store_buffer.sv:168:5
		req_port_o[2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1)))] = 1'b0;
		// Trace: core/store_buffer.sv:172:5
		if (commit_queue_q[(commit_read_pointer_q * ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 3 : 1 - (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2))) + ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? 0 : ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2)] && !stall_st_pending_i) begin
			// Trace: core/store_buffer.sv:173:7
			req_port_o[2 + ((dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[17102-:32] / 8) + (2 + (dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_dcache_req_i_t_CVA6Cfg[1124-:32] + 1)))] = 1'b1;
			// Trace: core/store_buffer.sv:174:7
			if (req_port_i[2 + (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[1124-:32] + (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[17102-:32] + (dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_dcache_req_o_t_CVA6Cfg[900-:32] - 1)))]) begin
				// Trace: core/store_buffer.sv:176:9
				commit_queue_n[(commit_read_pointer_q * ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 3 : 1 - (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2))) + ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? 0 : ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2)] = 1'b0;
				// Trace: core/store_buffer.sv:178:9
				commit_read_pointer_n = commit_read_pointer_q + 1'b1;
				// Trace: core/store_buffer.sv:179:9
				commit_status_cnt = commit_status_cnt - 1;
			end
		end
		if (commit_i) begin
			// Trace: core/store_buffer.sv:187:7
			commit_queue_n[((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? 0 : ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) + (commit_write_pointer_q * ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 3 : 1 - (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2)))+:((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 3 : 1 - (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2))] = speculative_queue_q[((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? 0 : ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) + (speculative_read_pointer_q * ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 3 : 1 - (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2)))+:((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 3 : 1 - (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2))];
			// Trace: core/store_buffer.sv:188:7
			commit_write_pointer_n = commit_write_pointer_n + 1'b1;
			// Trace: core/store_buffer.sv:189:7
			commit_status_cnt = commit_status_cnt + 1;
		end
		// Trace: core/store_buffer.sv:192:5
		commit_status_cnt_n = commit_status_cnt;
	end
	// Trace: core/store_buffer.sv:210:3
	always @(*) begin : sv2v_autoblock_2
		reg [0:1] _sv2v_jump;
		_sv2v_jump = 2'b00;
		begin : address_checker
			if (_sv2v_0)
				;
			// Trace: core/store_buffer.sv:211:5
			page_offset_matches_o = 1'b0;
			// Trace: core/store_buffer.sv:214:5
			begin : sv2v_autoblock_3
				// Trace: core/store_buffer.sv:214:10
				reg [31:0] i;
				// Trace: core/store_buffer.sv:214:10
				begin : sv2v_autoblock_4
					reg [31:0] _sv2v_value_on_break;
					for (i = 0; i < ariane_pkg_DEPTH_COMMIT; i = i + 1)
						if (_sv2v_jump < 2'b10) begin
							_sv2v_jump = 2'b00;
							// Trace: core/store_buffer.sv:216:7
							if ((page_offset_i[11:3] == commit_queue_q[((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? (i * ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 3 : 1 - (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2))) + ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12)) >= ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 4)) ? (CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12) : (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12)) + (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12)) >= ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 4)) ? (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12)) - ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 4))) + 1 : (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 4)) - ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12))) + 1)) - 1) : (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) - (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12)) >= ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 4)) ? (CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12) : (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12)) + (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12)) >= ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 4)) ? (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12)) - ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 4))) + 1 : (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 4)) - ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12))) + 1)) - 1)) : (((i * ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 3 : 1 - (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2))) + ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12)) >= ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 4)) ? (CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12) : (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12)) + (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12)) >= ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 4)) ? (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12)) - ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 4))) + 1 : (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 4)) - ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12))) + 1)) - 1) : (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) - (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12)) >= ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 4)) ? (CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12) : (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12)) + (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12)) >= ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 4)) ? (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12)) - ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 4))) + 1 : (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 4)) - ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12))) + 1)) - 1))) + (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12)) >= ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 4)) ? (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12)) - ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 4))) + 1 : (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 4)) - ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12))) + 1)) - 1)-:(((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12)) >= ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 4)) ? (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12)) - ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 4))) + 1 : (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 4)) - ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12))) + 1)]) && commit_queue_q[(i * ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 3 : 1 - (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2))) + ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? 0 : ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2)]) begin
								// Trace: core/store_buffer.sv:217:9
								page_offset_matches_o = 1'b1;
								// Trace: core/store_buffer.sv:218:9
								_sv2v_jump = 2'b10;
							end
							_sv2v_value_on_break = i;
						end
					if (!(_sv2v_jump < 2'b10))
						i = _sv2v_value_on_break;
					if (_sv2v_jump != 2'b11)
						_sv2v_jump = 2'b00;
				end
			end
			if (_sv2v_jump == 2'b00) begin
				begin : sv2v_autoblock_5
					// Trace: core/store_buffer.sv:222:10
					reg [31:0] i;
					// Trace: core/store_buffer.sv:222:10
					begin : sv2v_autoblock_6
						reg [31:0] _sv2v_value_on_break;
						for (i = 0; i < ariane_pkg_DEPTH_SPEC; i = i + 1)
							if (_sv2v_jump < 2'b10) begin
								_sv2v_jump = 2'b00;
								// Trace: core/store_buffer.sv:224:7
								if ((page_offset_i[11:3] == speculative_queue_q[((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? (i * ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 3 : 1 - (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2))) + ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12)) >= ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 4)) ? (CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12) : (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12)) + (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12)) >= ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 4)) ? (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12)) - ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 4))) + 1 : (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 4)) - ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12))) + 1)) - 1) : (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) - (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12)) >= ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 4)) ? (CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12) : (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12)) + (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12)) >= ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 4)) ? (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12)) - ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 4))) + 1 : (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 4)) - ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12))) + 1)) - 1)) : (((i * ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 3 : 1 - (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2))) + ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12)) >= ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 4)) ? (CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12) : (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12)) + (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12)) >= ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 4)) ? (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12)) - ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 4))) + 1 : (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 4)) - ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12))) + 1)) - 1) : (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) - (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12)) >= ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 4)) ? (CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12) : (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12)) + (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12)) >= ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 4)) ? (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12)) - ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 4))) + 1 : (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 4)) - ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12))) + 1)) - 1))) + (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12)) >= ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 4)) ? (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12)) - ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 4))) + 1 : (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 4)) - ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12))) + 1)) - 1)-:(((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12)) >= ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 4)) ? (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12)) - ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 4))) + 1 : (((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 4)) - ((CVA6Cfg[17038-:32] + (CVA6Cfg[17102-:32] + ((CVA6Cfg[17102-:32] / 8) + 2))) - (CVA6Cfg[17038-:32] - 12))) + 1)]) && speculative_queue_q[(i * ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 3 : 1 - (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2))) + ((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? 0 : ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2)]) begin
									// Trace: core/store_buffer.sv:225:9
									page_offset_matches_o = 1'b1;
									// Trace: core/store_buffer.sv:226:9
									_sv2v_jump = 2'b10;
								end
								_sv2v_value_on_break = i;
							end
						if (!(_sv2v_jump < 2'b10))
							i = _sv2v_value_on_break;
						if (_sv2v_jump != 2'b11)
							_sv2v_jump = 2'b00;
					end
				end
				if (_sv2v_jump == 2'b00) begin
					if ((page_offset_i[11:3] == paddr_i[11:3]) && valid_without_flush_i)
						// Trace: core/store_buffer.sv:231:7
						page_offset_matches_o = 1'b1;
				end
			end
		end
	end
	// Trace: core/store_buffer.sv:237:3
	function automatic [((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 3 : 1 - (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2)) - 1:0] sv2v_cast_6EC44;
		input reg [((((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2) >= 0 ? ((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 3 : 1 - (((CVA6Cfg[17038-:32] + CVA6Cfg[17102-:32]) + (CVA6Cfg[17102-:32] / 8)) + 2)) - 1:0] inp;
		sv2v_cast_6EC44 = inp;
	endfunction
	always @(posedge clk_i or negedge rst_ni) begin : p_spec
		// Trace: core/store_buffer.sv:238:5
		if (~rst_ni) begin
			// Trace: core/store_buffer.sv:239:7
			speculative_queue_q <= {ariane_pkg_DEPTH_SPEC {sv2v_cast_6EC44(0)}};
			// Trace: core/store_buffer.sv:240:7
			speculative_read_pointer_q <= 1'sb0;
			// Trace: core/store_buffer.sv:241:7
			speculative_write_pointer_q <= 1'sb0;
			// Trace: core/store_buffer.sv:242:7
			speculative_status_cnt_q <= 1'sb0;
		end
		else begin
			// Trace: core/store_buffer.sv:244:7
			speculative_queue_q <= speculative_queue_n;
			// Trace: core/store_buffer.sv:245:7
			speculative_read_pointer_q <= speculative_read_pointer_n;
			// Trace: core/store_buffer.sv:246:7
			speculative_write_pointer_q <= speculative_write_pointer_n;
			// Trace: core/store_buffer.sv:247:7
			speculative_status_cnt_q <= speculative_status_cnt_n;
		end
	end
	// Trace: core/store_buffer.sv:252:3
	always @(posedge clk_i or negedge rst_ni) begin : p_commit
		// Trace: core/store_buffer.sv:253:5
		if (~rst_ni) begin
			// Trace: core/store_buffer.sv:254:7
			commit_queue_q <= {ariane_pkg_DEPTH_COMMIT {sv2v_cast_6EC44(0)}};
			// Trace: core/store_buffer.sv:255:7
			commit_read_pointer_q <= 1'sb0;
			// Trace: core/store_buffer.sv:256:7
			commit_write_pointer_q <= 1'sb0;
			// Trace: core/store_buffer.sv:257:7
			commit_status_cnt_q <= 1'sb0;
		end
		else begin
			// Trace: core/store_buffer.sv:259:7
			commit_queue_q <= commit_queue_n;
			// Trace: core/store_buffer.sv:260:7
			commit_read_pointer_q <= commit_read_pointer_n;
			// Trace: core/store_buffer.sv:261:7
			commit_write_pointer_q <= commit_write_pointer_n;
			// Trace: core/store_buffer.sv:262:7
			commit_status_cnt_q <= commit_status_cnt_n;
		end
	end
	// Trace: core/store_buffer.sv:273:3
	// removed an assertion item
	// commit_and_flush : assert property (@(posedge clk_i) 
	// 	(rst_ni && flush_i |-> !commit_i)
	// ) else begin
	// 	// Trace: core/store_buffer.sv:275:8
	// 	$error("[Commit Queue] You are trying to commit and flush in the same cycle");
	// end
	// Trace: core/store_buffer.sv:277:3
	// removed an assertion item
	// speculative_buffer_overflow : assert property (@(posedge clk_i) 
	// 	(rst_ni && (speculative_status_cnt_q == ariane_pkg_DEPTH_SPEC) |-> !valid_i)
	// ) else begin
	// 	// Trace: core/store_buffer.sv:280:5
	// 	$error("[Speculative Queue] You are trying to push new data although the buffer is not ready");
	// end
	// Trace: core/store_buffer.sv:282:3
	// removed an assertion item
	// speculative_buffer_underflow : assert property (@(posedge clk_i) 
	// 	(rst_ni && (speculative_status_cnt_q == 0) |-> !commit_i)
	// ) else begin
	// 	// Trace: core/store_buffer.sv:284:8
	// 	$error("[Speculative Queue] You are committing although there are no stores to commit");
	// end
	// Trace: core/store_buffer.sv:286:3
	// removed an assertion item
	// commit_buffer_overflow : assert property (@(posedge clk_i) 
	// 	(rst_ni && (commit_status_cnt_q == ariane_pkg_DEPTH_COMMIT) |-> !commit_i)
	// ) else begin
	// 	// Trace: core/store_buffer.sv:288:8
	// 	$error("[Commit Queue] You are trying to commit a store although the buffer is full");
	// end
	initial _sv2v_0 = 0;
endmodule
