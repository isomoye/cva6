// removed module with interface ports: axi2mem
